module BTB(input clk, input reset,
    input  io_req_valid,
    input [42:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output io_resp_bits_mask,
    output io_resp_bits_bridx,
    output[42:0] io_resp_bits_target,
    output[5:0] io_resp_bits_entry,
    output[6:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_btb_update_valid,
    input  io_btb_update_bits_prediction_valid,
    input  io_btb_update_bits_prediction_bits_taken,
    input  io_btb_update_bits_prediction_bits_mask,
    input  io_btb_update_bits_prediction_bits_bridx,
    input [42:0] io_btb_update_bits_prediction_bits_target,
    input [5:0] io_btb_update_bits_prediction_bits_entry,
    input [6:0] io_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_btb_update_bits_pc,
    input [42:0] io_btb_update_bits_target,
    input  io_btb_update_bits_taken,
    input  io_btb_update_bits_isJump,
    input  io_btb_update_bits_isReturn,
    input [42:0] io_btb_update_bits_br_pc,
    input  io_bht_update_valid,
    input  io_bht_update_bits_prediction_valid,
    input  io_bht_update_bits_prediction_bits_taken,
    input  io_bht_update_bits_prediction_bits_mask,
    input  io_bht_update_bits_prediction_bits_bridx,
    input [42:0] io_bht_update_bits_prediction_bits_target,
    input [5:0] io_bht_update_bits_prediction_bits_entry,
    input [6:0] io_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_bht_update_bits_prediction_bits_bht_value,
    input [42:0] io_bht_update_bits_pc,
    input  io_bht_update_bits_taken,
    input  io_bht_update_bits_mispredict,
    input  io_ras_update_valid,
    input  io_ras_update_bits_isCall,
    input  io_ras_update_bits_isReturn,
    input [42:0] io_ras_update_bits_returnAddr,
    input  io_ras_update_bits_prediction_valid,
    input  io_ras_update_bits_prediction_bits_taken,
    input  io_ras_update_bits_prediction_bits_mask,
    input  io_ras_update_bits_prediction_bits_bridx,
    input [42:0] io_ras_update_bits_prediction_bits_target,
    input [5:0] io_ras_update_bits_prediction_bits_entry,
    input [6:0] io_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_ras_update_bits_prediction_bits_bht_value,
    input  io_invalidate
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg [42:0] R4;
  wire[42:0] T5;
  wire T6;
  reg  R7;
  wire T1579;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10 [127:0];
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[6:0] T24;
  reg [6:0] R25;
  wire[6:0] T26;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[5:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[61:0] T34;
  reg [61:0] isJump;
  wire[61:0] T1580;
  wire[63:0] T35;
  wire[63:0] T1581;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T1582;
  wire[61:0] T39;
  wire[63:0] T40;
  wire[5:0] T41;
  reg [5:0] R42;
  wire[5:0] T1583;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire T46;
  wire T47;
  wire T48;
  reg [5:0] R49;
  wire[5:0] T50;
  reg  updateHit;
  wire T51;
  wire[63:0] T1584;
  wire T52;
  wire T53;
  reg  R54;
  wire T55;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T1585;
  wire[61:0] hits;
  wire[61:0] T58;
  wire[61:0] T59;
  wire[30:0] T60;
  wire[15:0] T61;
  wire[7:0] T62;
  wire[3:0] T63;
  wire[1:0] T64;
  wire T65;
  wire[5:0] T66;
  wire[5:0] pageHit;
  reg [5:0] pageValid;
  wire[5:0] T1586;
  wire[7:0] T1587;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T1588;
  wire[7:0] T69;
  wire[7:0] pageReplEn;
  wire[7:0] tgtPageReplEn;
  wire[7:0] tgtPageRepl;
  wire[7:0] T1589;
  wire[5:0] T70;
  wire[5:0] T1590;
  wire T71;
  wire[5:0] T72;
  wire[4:0] T73;
  wire[7:0] idxPageUpdateOH;
  wire[7:0] idxPageRepl;
  wire[7:0] T74;
  reg [2:0] R75;
  wire[2:0] T1591;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire[7:0] T1592;
  wire[5:0] updatePageHit;
  wire[5:0] T81;
  wire[5:0] T82;
  wire[2:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[29:0] T86;
  reg [42:0] R87;
  wire[42:0] T88;
  wire[29:0] T89;
  reg [29:0] pages [5:0];
  wire[29:0] T90;
  wire[29:0] T91;
  wire[29:0] T92;
  wire[29:0] T93;
  wire T94;
  wire[7:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[29:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire[29:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[29:0] T108;
  wire[29:0] T109;
  wire[29:0] T110;
  wire[29:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[29:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire[29:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[29:0] T125;
  wire T126;
  wire[29:0] T127;
  wire[2:0] T128;
  wire[1:0] T129;
  wire T130;
  wire[29:0] T131;
  wire T132;
  wire[29:0] T133;
  wire T134;
  wire[29:0] T135;
  wire useUpdatePageHit;
  wire samePage;
  wire[29:0] T136;
  wire[29:0] T137;
  wire doTgtPageRepl;
  wire T138;
  wire usePageHit;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[7:0] T1593;
  wire T141;
  wire[7:0] idxPageReplEn;
  wire[7:0] T1594;
  wire T142;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  wire T147;
  wire[29:0] T148;
  wire[29:0] T149;
  wire T150;
  wire[29:0] T151;
  wire T152;
  wire[29:0] T153;
  wire[2:0] T154;
  wire[1:0] T155;
  wire T156;
  wire[29:0] T157;
  wire T158;
  wire[29:0] T159;
  wire T160;
  wire[29:0] T161;
  wire[5:0] idxPagesOH_0;
  wire[7:0] T162;
  wire[2:0] T163;
  reg [2:0] idxPages [61:0];
  wire[2:0] T164;
  wire[2:0] T1595;
  wire[1:0] T1596;
  wire T1597;
  wire[1:0] T1598;
  wire[1:0] T1599;
  wire[3:0] T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[1:0] T1603;
  wire T1604;
  wire T1605;
  wire T165;
  wire T166;
  wire T167;
  wire[5:0] T168;
  wire[5:0] idxPagesOH_1;
  wire[7:0] T169;
  wire[2:0] T170;
  wire[1:0] T171;
  wire T172;
  wire[5:0] T173;
  wire[5:0] idxPagesOH_2;
  wire[7:0] T174;
  wire[2:0] T175;
  wire T176;
  wire[5:0] T177;
  wire[5:0] idxPagesOH_3;
  wire[7:0] T178;
  wire[2:0] T179;
  wire[3:0] T180;
  wire[1:0] T181;
  wire T182;
  wire[5:0] T183;
  wire[5:0] idxPagesOH_4;
  wire[7:0] T184;
  wire[2:0] T185;
  wire T186;
  wire[5:0] T187;
  wire[5:0] idxPagesOH_5;
  wire[7:0] T188;
  wire[2:0] T189;
  wire[1:0] T190;
  wire T191;
  wire[5:0] T192;
  wire[5:0] idxPagesOH_6;
  wire[7:0] T193;
  wire[2:0] T194;
  wire T195;
  wire[5:0] T196;
  wire[5:0] idxPagesOH_7;
  wire[7:0] T197;
  wire[2:0] T198;
  wire[7:0] T199;
  wire[3:0] T200;
  wire[1:0] T201;
  wire T202;
  wire[5:0] T203;
  wire[5:0] idxPagesOH_8;
  wire[7:0] T204;
  wire[2:0] T205;
  wire T206;
  wire[5:0] T207;
  wire[5:0] idxPagesOH_9;
  wire[7:0] T208;
  wire[2:0] T209;
  wire[1:0] T210;
  wire T211;
  wire[5:0] T212;
  wire[5:0] idxPagesOH_10;
  wire[7:0] T213;
  wire[2:0] T214;
  wire T215;
  wire[5:0] T216;
  wire[5:0] idxPagesOH_11;
  wire[7:0] T217;
  wire[2:0] T218;
  wire[3:0] T219;
  wire[1:0] T220;
  wire T221;
  wire[5:0] T222;
  wire[5:0] idxPagesOH_12;
  wire[7:0] T223;
  wire[2:0] T224;
  wire T225;
  wire[5:0] T226;
  wire[5:0] idxPagesOH_13;
  wire[7:0] T227;
  wire[2:0] T228;
  wire[1:0] T229;
  wire T230;
  wire[5:0] T231;
  wire[5:0] idxPagesOH_14;
  wire[7:0] T232;
  wire[2:0] T233;
  wire T234;
  wire[5:0] T235;
  wire[5:0] idxPagesOH_15;
  wire[7:0] T236;
  wire[2:0] T237;
  wire[14:0] T238;
  wire[7:0] T239;
  wire[3:0] T240;
  wire[1:0] T241;
  wire T242;
  wire[5:0] T243;
  wire[5:0] idxPagesOH_16;
  wire[7:0] T244;
  wire[2:0] T245;
  wire T246;
  wire[5:0] T247;
  wire[5:0] idxPagesOH_17;
  wire[7:0] T248;
  wire[2:0] T249;
  wire[1:0] T250;
  wire T251;
  wire[5:0] T252;
  wire[5:0] idxPagesOH_18;
  wire[7:0] T253;
  wire[2:0] T254;
  wire T255;
  wire[5:0] T256;
  wire[5:0] idxPagesOH_19;
  wire[7:0] T257;
  wire[2:0] T258;
  wire[3:0] T259;
  wire[1:0] T260;
  wire T261;
  wire[5:0] T262;
  wire[5:0] idxPagesOH_20;
  wire[7:0] T263;
  wire[2:0] T264;
  wire T265;
  wire[5:0] T266;
  wire[5:0] idxPagesOH_21;
  wire[7:0] T267;
  wire[2:0] T268;
  wire[1:0] T269;
  wire T270;
  wire[5:0] T271;
  wire[5:0] idxPagesOH_22;
  wire[7:0] T272;
  wire[2:0] T273;
  wire T274;
  wire[5:0] T275;
  wire[5:0] idxPagesOH_23;
  wire[7:0] T276;
  wire[2:0] T277;
  wire[6:0] T278;
  wire[3:0] T279;
  wire[1:0] T280;
  wire T281;
  wire[5:0] T282;
  wire[5:0] idxPagesOH_24;
  wire[7:0] T283;
  wire[2:0] T284;
  wire T285;
  wire[5:0] T286;
  wire[5:0] idxPagesOH_25;
  wire[7:0] T287;
  wire[2:0] T288;
  wire[1:0] T289;
  wire T290;
  wire[5:0] T291;
  wire[5:0] idxPagesOH_26;
  wire[7:0] T292;
  wire[2:0] T293;
  wire T294;
  wire[5:0] T295;
  wire[5:0] idxPagesOH_27;
  wire[7:0] T296;
  wire[2:0] T297;
  wire[2:0] T298;
  wire[1:0] T299;
  wire T300;
  wire[5:0] T301;
  wire[5:0] idxPagesOH_28;
  wire[7:0] T302;
  wire[2:0] T303;
  wire T304;
  wire[5:0] T305;
  wire[5:0] idxPagesOH_29;
  wire[7:0] T306;
  wire[2:0] T307;
  wire T308;
  wire[5:0] T309;
  wire[5:0] idxPagesOH_30;
  wire[7:0] T310;
  wire[2:0] T311;
  wire[30:0] T312;
  wire[15:0] T313;
  wire[7:0] T314;
  wire[3:0] T315;
  wire[1:0] T316;
  wire T317;
  wire[5:0] T318;
  wire[5:0] idxPagesOH_31;
  wire[7:0] T319;
  wire[2:0] T320;
  wire T321;
  wire[5:0] T322;
  wire[5:0] idxPagesOH_32;
  wire[7:0] T323;
  wire[2:0] T324;
  wire[1:0] T325;
  wire T326;
  wire[5:0] T327;
  wire[5:0] idxPagesOH_33;
  wire[7:0] T328;
  wire[2:0] T329;
  wire T330;
  wire[5:0] T331;
  wire[5:0] idxPagesOH_34;
  wire[7:0] T332;
  wire[2:0] T333;
  wire[3:0] T334;
  wire[1:0] T335;
  wire T336;
  wire[5:0] T337;
  wire[5:0] idxPagesOH_35;
  wire[7:0] T338;
  wire[2:0] T339;
  wire T340;
  wire[5:0] T341;
  wire[5:0] idxPagesOH_36;
  wire[7:0] T342;
  wire[2:0] T343;
  wire[1:0] T344;
  wire T345;
  wire[5:0] T346;
  wire[5:0] idxPagesOH_37;
  wire[7:0] T347;
  wire[2:0] T348;
  wire T349;
  wire[5:0] T350;
  wire[5:0] idxPagesOH_38;
  wire[7:0] T351;
  wire[2:0] T352;
  wire[7:0] T353;
  wire[3:0] T354;
  wire[1:0] T355;
  wire T356;
  wire[5:0] T357;
  wire[5:0] idxPagesOH_39;
  wire[7:0] T358;
  wire[2:0] T359;
  wire T360;
  wire[5:0] T361;
  wire[5:0] idxPagesOH_40;
  wire[7:0] T362;
  wire[2:0] T363;
  wire[1:0] T364;
  wire T365;
  wire[5:0] T366;
  wire[5:0] idxPagesOH_41;
  wire[7:0] T367;
  wire[2:0] T368;
  wire T369;
  wire[5:0] T370;
  wire[5:0] idxPagesOH_42;
  wire[7:0] T371;
  wire[2:0] T372;
  wire[3:0] T373;
  wire[1:0] T374;
  wire T375;
  wire[5:0] T376;
  wire[5:0] idxPagesOH_43;
  wire[7:0] T377;
  wire[2:0] T378;
  wire T379;
  wire[5:0] T380;
  wire[5:0] idxPagesOH_44;
  wire[7:0] T381;
  wire[2:0] T382;
  wire[1:0] T383;
  wire T384;
  wire[5:0] T385;
  wire[5:0] idxPagesOH_45;
  wire[7:0] T386;
  wire[2:0] T387;
  wire T388;
  wire[5:0] T389;
  wire[5:0] idxPagesOH_46;
  wire[7:0] T390;
  wire[2:0] T391;
  wire[14:0] T392;
  wire[7:0] T393;
  wire[3:0] T394;
  wire[1:0] T395;
  wire T396;
  wire[5:0] T397;
  wire[5:0] idxPagesOH_47;
  wire[7:0] T398;
  wire[2:0] T399;
  wire T400;
  wire[5:0] T401;
  wire[5:0] idxPagesOH_48;
  wire[7:0] T402;
  wire[2:0] T403;
  wire[1:0] T404;
  wire T405;
  wire[5:0] T406;
  wire[5:0] idxPagesOH_49;
  wire[7:0] T407;
  wire[2:0] T408;
  wire T409;
  wire[5:0] T410;
  wire[5:0] idxPagesOH_50;
  wire[7:0] T411;
  wire[2:0] T412;
  wire[3:0] T413;
  wire[1:0] T414;
  wire T415;
  wire[5:0] T416;
  wire[5:0] idxPagesOH_51;
  wire[7:0] T417;
  wire[2:0] T418;
  wire T419;
  wire[5:0] T420;
  wire[5:0] idxPagesOH_52;
  wire[7:0] T421;
  wire[2:0] T422;
  wire[1:0] T423;
  wire T424;
  wire[5:0] T425;
  wire[5:0] idxPagesOH_53;
  wire[7:0] T426;
  wire[2:0] T427;
  wire T428;
  wire[5:0] T429;
  wire[5:0] idxPagesOH_54;
  wire[7:0] T430;
  wire[2:0] T431;
  wire[6:0] T432;
  wire[3:0] T433;
  wire[1:0] T434;
  wire T435;
  wire[5:0] T436;
  wire[5:0] idxPagesOH_55;
  wire[7:0] T437;
  wire[2:0] T438;
  wire T439;
  wire[5:0] T440;
  wire[5:0] idxPagesOH_56;
  wire[7:0] T441;
  wire[2:0] T442;
  wire[1:0] T443;
  wire T444;
  wire[5:0] T445;
  wire[5:0] idxPagesOH_57;
  wire[7:0] T446;
  wire[2:0] T447;
  wire T448;
  wire[5:0] T449;
  wire[5:0] idxPagesOH_58;
  wire[7:0] T450;
  wire[2:0] T451;
  wire[2:0] T452;
  wire[1:0] T453;
  wire T454;
  wire[5:0] T455;
  wire[5:0] idxPagesOH_59;
  wire[7:0] T456;
  wire[2:0] T457;
  wire T458;
  wire[5:0] T459;
  wire[5:0] idxPagesOH_60;
  wire[7:0] T460;
  wire[2:0] T461;
  wire T462;
  wire[5:0] T463;
  wire[5:0] idxPagesOH_61;
  wire[7:0] T464;
  wire[2:0] T465;
  wire[61:0] T466;
  wire[61:0] T467;
  wire[61:0] T468;
  wire[30:0] T469;
  wire[15:0] T470;
  wire[7:0] T471;
  wire[3:0] T472;
  wire[1:0] T473;
  wire T474;
  wire[12:0] T475;
  wire[12:0] T476;
  reg [12:0] idxs [61:0];
  wire[12:0] T477;
  wire[12:0] T1606;
  wire T478;
  wire T479;
  wire T480;
  wire[12:0] T481;
  wire[1:0] T482;
  wire T483;
  wire[12:0] T484;
  wire T485;
  wire[12:0] T486;
  wire[3:0] T487;
  wire[1:0] T488;
  wire T489;
  wire[12:0] T490;
  wire T491;
  wire[12:0] T492;
  wire[1:0] T493;
  wire T494;
  wire[12:0] T495;
  wire T496;
  wire[12:0] T497;
  wire[7:0] T498;
  wire[3:0] T499;
  wire[1:0] T500;
  wire T501;
  wire[12:0] T502;
  wire T503;
  wire[12:0] T504;
  wire[1:0] T505;
  wire T506;
  wire[12:0] T507;
  wire T508;
  wire[12:0] T509;
  wire[3:0] T510;
  wire[1:0] T511;
  wire T512;
  wire[12:0] T513;
  wire T514;
  wire[12:0] T515;
  wire[1:0] T516;
  wire T517;
  wire[12:0] T518;
  wire T519;
  wire[12:0] T520;
  wire[14:0] T521;
  wire[7:0] T522;
  wire[3:0] T523;
  wire[1:0] T524;
  wire T525;
  wire[12:0] T526;
  wire T527;
  wire[12:0] T528;
  wire[1:0] T529;
  wire T530;
  wire[12:0] T531;
  wire T532;
  wire[12:0] T533;
  wire[3:0] T534;
  wire[1:0] T535;
  wire T536;
  wire[12:0] T537;
  wire T538;
  wire[12:0] T539;
  wire[1:0] T540;
  wire T541;
  wire[12:0] T542;
  wire T543;
  wire[12:0] T544;
  wire[6:0] T545;
  wire[3:0] T546;
  wire[1:0] T547;
  wire T548;
  wire[12:0] T549;
  wire T550;
  wire[12:0] T551;
  wire[1:0] T552;
  wire T553;
  wire[12:0] T554;
  wire T555;
  wire[12:0] T556;
  wire[2:0] T557;
  wire[1:0] T558;
  wire T559;
  wire[12:0] T560;
  wire T561;
  wire[12:0] T562;
  wire T563;
  wire[12:0] T564;
  wire[30:0] T565;
  wire[15:0] T566;
  wire[7:0] T567;
  wire[3:0] T568;
  wire[1:0] T569;
  wire T570;
  wire[12:0] T571;
  wire T572;
  wire[12:0] T573;
  wire[1:0] T574;
  wire T575;
  wire[12:0] T576;
  wire T577;
  wire[12:0] T578;
  wire[3:0] T579;
  wire[1:0] T580;
  wire T581;
  wire[12:0] T582;
  wire T583;
  wire[12:0] T584;
  wire[1:0] T585;
  wire T586;
  wire[12:0] T587;
  wire T588;
  wire[12:0] T589;
  wire[7:0] T590;
  wire[3:0] T591;
  wire[1:0] T592;
  wire T593;
  wire[12:0] T594;
  wire T595;
  wire[12:0] T596;
  wire[1:0] T597;
  wire T598;
  wire[12:0] T599;
  wire T600;
  wire[12:0] T601;
  wire[3:0] T602;
  wire[1:0] T603;
  wire T604;
  wire[12:0] T605;
  wire T606;
  wire[12:0] T607;
  wire[1:0] T608;
  wire T609;
  wire[12:0] T610;
  wire T611;
  wire[12:0] T612;
  wire[14:0] T613;
  wire[7:0] T614;
  wire[3:0] T615;
  wire[1:0] T616;
  wire T617;
  wire[12:0] T618;
  wire T619;
  wire[12:0] T620;
  wire[1:0] T621;
  wire T622;
  wire[12:0] T623;
  wire T624;
  wire[12:0] T625;
  wire[3:0] T626;
  wire[1:0] T627;
  wire T628;
  wire[12:0] T629;
  wire T630;
  wire[12:0] T631;
  wire[1:0] T632;
  wire T633;
  wire[12:0] T634;
  wire T635;
  wire[12:0] T636;
  wire[6:0] T637;
  wire[3:0] T638;
  wire[1:0] T639;
  wire T640;
  wire[12:0] T641;
  wire T642;
  wire[12:0] T643;
  wire[1:0] T644;
  wire T645;
  wire[12:0] T646;
  wire T647;
  wire[12:0] T648;
  wire[2:0] T649;
  wire[1:0] T650;
  wire T651;
  wire[12:0] T652;
  wire T653;
  wire[12:0] T654;
  wire T655;
  wire[12:0] T656;
  reg [61:0] idxValid;
  wire[61:0] T1607;
  wire[63:0] T1608;
  wire[63:0] T657;
  wire[63:0] T658;
  wire[63:0] T1609;
  wire[61:0] T659;
  wire[61:0] T660;
  wire[61:0] T661;
  wire[61:0] T662;
  wire[61:0] T663;
  wire[30:0] T664;
  wire[15:0] T665;
  wire[7:0] T666;
  wire[3:0] T667;
  wire[1:0] T668;
  wire T669;
  wire[7:0] T670;
  wire[7:0] T1610;
  wire[5:0] T671;
  wire[5:0] tgtPagesOH_0;
  wire[7:0] T672;
  wire[2:0] T673;
  reg [2:0] tgtPages [61:0];
  wire[2:0] T674;
  wire[2:0] T1611;
  wire[1:0] T1612;
  wire T1613;
  wire[1:0] T1614;
  wire[1:0] T1615;
  wire[3:0] T1616;
  wire[3:0] T1617;
  wire[7:0] T675;
  wire[7:0] T1618;
  wire[3:0] T1619;
  wire[1:0] T1620;
  wire T1621;
  wire T1622;
  wire T676;
  wire T677;
  wire T678;
  wire[7:0] T679;
  wire[7:0] T1623;
  wire[5:0] T680;
  wire[5:0] tgtPagesOH_1;
  wire[7:0] T681;
  wire[2:0] T682;
  wire[1:0] T683;
  wire T684;
  wire[7:0] T685;
  wire[7:0] T1624;
  wire[5:0] T686;
  wire[5:0] tgtPagesOH_2;
  wire[7:0] T687;
  wire[2:0] T688;
  wire T689;
  wire[7:0] T690;
  wire[7:0] T1625;
  wire[5:0] T691;
  wire[5:0] tgtPagesOH_3;
  wire[7:0] T692;
  wire[2:0] T693;
  wire[3:0] T694;
  wire[1:0] T695;
  wire T696;
  wire[7:0] T697;
  wire[7:0] T1626;
  wire[5:0] T698;
  wire[5:0] tgtPagesOH_4;
  wire[7:0] T699;
  wire[2:0] T700;
  wire T701;
  wire[7:0] T702;
  wire[7:0] T1627;
  wire[5:0] T703;
  wire[5:0] tgtPagesOH_5;
  wire[7:0] T704;
  wire[2:0] T705;
  wire[1:0] T706;
  wire T707;
  wire[7:0] T708;
  wire[7:0] T1628;
  wire[5:0] T709;
  wire[5:0] tgtPagesOH_6;
  wire[7:0] T710;
  wire[2:0] T711;
  wire T712;
  wire[7:0] T713;
  wire[7:0] T1629;
  wire[5:0] T714;
  wire[5:0] tgtPagesOH_7;
  wire[7:0] T715;
  wire[2:0] T716;
  wire[7:0] T717;
  wire[3:0] T718;
  wire[1:0] T719;
  wire T720;
  wire[7:0] T721;
  wire[7:0] T1630;
  wire[5:0] T722;
  wire[5:0] tgtPagesOH_8;
  wire[7:0] T723;
  wire[2:0] T724;
  wire T725;
  wire[7:0] T726;
  wire[7:0] T1631;
  wire[5:0] T727;
  wire[5:0] tgtPagesOH_9;
  wire[7:0] T728;
  wire[2:0] T729;
  wire[1:0] T730;
  wire T731;
  wire[7:0] T732;
  wire[7:0] T1632;
  wire[5:0] T733;
  wire[5:0] tgtPagesOH_10;
  wire[7:0] T734;
  wire[2:0] T735;
  wire T736;
  wire[7:0] T737;
  wire[7:0] T1633;
  wire[5:0] T738;
  wire[5:0] tgtPagesOH_11;
  wire[7:0] T739;
  wire[2:0] T740;
  wire[3:0] T741;
  wire[1:0] T742;
  wire T743;
  wire[7:0] T744;
  wire[7:0] T1634;
  wire[5:0] T745;
  wire[5:0] tgtPagesOH_12;
  wire[7:0] T746;
  wire[2:0] T747;
  wire T748;
  wire[7:0] T749;
  wire[7:0] T1635;
  wire[5:0] T750;
  wire[5:0] tgtPagesOH_13;
  wire[7:0] T751;
  wire[2:0] T752;
  wire[1:0] T753;
  wire T754;
  wire[7:0] T755;
  wire[7:0] T1636;
  wire[5:0] T756;
  wire[5:0] tgtPagesOH_14;
  wire[7:0] T757;
  wire[2:0] T758;
  wire T759;
  wire[7:0] T760;
  wire[7:0] T1637;
  wire[5:0] T761;
  wire[5:0] tgtPagesOH_15;
  wire[7:0] T762;
  wire[2:0] T763;
  wire[14:0] T764;
  wire[7:0] T765;
  wire[3:0] T766;
  wire[1:0] T767;
  wire T768;
  wire[7:0] T769;
  wire[7:0] T1638;
  wire[5:0] T770;
  wire[5:0] tgtPagesOH_16;
  wire[7:0] T771;
  wire[2:0] T772;
  wire T773;
  wire[7:0] T774;
  wire[7:0] T1639;
  wire[5:0] T775;
  wire[5:0] tgtPagesOH_17;
  wire[7:0] T776;
  wire[2:0] T777;
  wire[1:0] T778;
  wire T779;
  wire[7:0] T780;
  wire[7:0] T1640;
  wire[5:0] T781;
  wire[5:0] tgtPagesOH_18;
  wire[7:0] T782;
  wire[2:0] T783;
  wire T784;
  wire[7:0] T785;
  wire[7:0] T1641;
  wire[5:0] T786;
  wire[5:0] tgtPagesOH_19;
  wire[7:0] T787;
  wire[2:0] T788;
  wire[3:0] T789;
  wire[1:0] T790;
  wire T791;
  wire[7:0] T792;
  wire[7:0] T1642;
  wire[5:0] T793;
  wire[5:0] tgtPagesOH_20;
  wire[7:0] T794;
  wire[2:0] T795;
  wire T796;
  wire[7:0] T797;
  wire[7:0] T1643;
  wire[5:0] T798;
  wire[5:0] tgtPagesOH_21;
  wire[7:0] T799;
  wire[2:0] T800;
  wire[1:0] T801;
  wire T802;
  wire[7:0] T803;
  wire[7:0] T1644;
  wire[5:0] T804;
  wire[5:0] tgtPagesOH_22;
  wire[7:0] T805;
  wire[2:0] T806;
  wire T807;
  wire[7:0] T808;
  wire[7:0] T1645;
  wire[5:0] T809;
  wire[5:0] tgtPagesOH_23;
  wire[7:0] T810;
  wire[2:0] T811;
  wire[6:0] T812;
  wire[3:0] T813;
  wire[1:0] T814;
  wire T815;
  wire[7:0] T816;
  wire[7:0] T1646;
  wire[5:0] T817;
  wire[5:0] tgtPagesOH_24;
  wire[7:0] T818;
  wire[2:0] T819;
  wire T820;
  wire[7:0] T821;
  wire[7:0] T1647;
  wire[5:0] T822;
  wire[5:0] tgtPagesOH_25;
  wire[7:0] T823;
  wire[2:0] T824;
  wire[1:0] T825;
  wire T826;
  wire[7:0] T827;
  wire[7:0] T1648;
  wire[5:0] T828;
  wire[5:0] tgtPagesOH_26;
  wire[7:0] T829;
  wire[2:0] T830;
  wire T831;
  wire[7:0] T832;
  wire[7:0] T1649;
  wire[5:0] T833;
  wire[5:0] tgtPagesOH_27;
  wire[7:0] T834;
  wire[2:0] T835;
  wire[2:0] T836;
  wire[1:0] T837;
  wire T838;
  wire[7:0] T839;
  wire[7:0] T1650;
  wire[5:0] T840;
  wire[5:0] tgtPagesOH_28;
  wire[7:0] T841;
  wire[2:0] T842;
  wire T843;
  wire[7:0] T844;
  wire[7:0] T1651;
  wire[5:0] T845;
  wire[5:0] tgtPagesOH_29;
  wire[7:0] T846;
  wire[2:0] T847;
  wire T848;
  wire[7:0] T849;
  wire[7:0] T1652;
  wire[5:0] T850;
  wire[5:0] tgtPagesOH_30;
  wire[7:0] T851;
  wire[2:0] T852;
  wire[30:0] T853;
  wire[15:0] T854;
  wire[7:0] T855;
  wire[3:0] T856;
  wire[1:0] T857;
  wire T858;
  wire[7:0] T859;
  wire[7:0] T1653;
  wire[5:0] T860;
  wire[5:0] tgtPagesOH_31;
  wire[7:0] T861;
  wire[2:0] T862;
  wire T863;
  wire[7:0] T864;
  wire[7:0] T1654;
  wire[5:0] T865;
  wire[5:0] tgtPagesOH_32;
  wire[7:0] T866;
  wire[2:0] T867;
  wire[1:0] T868;
  wire T869;
  wire[7:0] T870;
  wire[7:0] T1655;
  wire[5:0] T871;
  wire[5:0] tgtPagesOH_33;
  wire[7:0] T872;
  wire[2:0] T873;
  wire T874;
  wire[7:0] T875;
  wire[7:0] T1656;
  wire[5:0] T876;
  wire[5:0] tgtPagesOH_34;
  wire[7:0] T877;
  wire[2:0] T878;
  wire[3:0] T879;
  wire[1:0] T880;
  wire T881;
  wire[7:0] T882;
  wire[7:0] T1657;
  wire[5:0] T883;
  wire[5:0] tgtPagesOH_35;
  wire[7:0] T884;
  wire[2:0] T885;
  wire T886;
  wire[7:0] T887;
  wire[7:0] T1658;
  wire[5:0] T888;
  wire[5:0] tgtPagesOH_36;
  wire[7:0] T889;
  wire[2:0] T890;
  wire[1:0] T891;
  wire T892;
  wire[7:0] T893;
  wire[7:0] T1659;
  wire[5:0] T894;
  wire[5:0] tgtPagesOH_37;
  wire[7:0] T895;
  wire[2:0] T896;
  wire T897;
  wire[7:0] T898;
  wire[7:0] T1660;
  wire[5:0] T899;
  wire[5:0] tgtPagesOH_38;
  wire[7:0] T900;
  wire[2:0] T901;
  wire[7:0] T902;
  wire[3:0] T903;
  wire[1:0] T904;
  wire T905;
  wire[7:0] T906;
  wire[7:0] T1661;
  wire[5:0] T907;
  wire[5:0] tgtPagesOH_39;
  wire[7:0] T908;
  wire[2:0] T909;
  wire T910;
  wire[7:0] T911;
  wire[7:0] T1662;
  wire[5:0] T912;
  wire[5:0] tgtPagesOH_40;
  wire[7:0] T913;
  wire[2:0] T914;
  wire[1:0] T915;
  wire T916;
  wire[7:0] T917;
  wire[7:0] T1663;
  wire[5:0] T918;
  wire[5:0] tgtPagesOH_41;
  wire[7:0] T919;
  wire[2:0] T920;
  wire T921;
  wire[7:0] T922;
  wire[7:0] T1664;
  wire[5:0] T923;
  wire[5:0] tgtPagesOH_42;
  wire[7:0] T924;
  wire[2:0] T925;
  wire[3:0] T926;
  wire[1:0] T927;
  wire T928;
  wire[7:0] T929;
  wire[7:0] T1665;
  wire[5:0] T930;
  wire[5:0] tgtPagesOH_43;
  wire[7:0] T931;
  wire[2:0] T932;
  wire T933;
  wire[7:0] T934;
  wire[7:0] T1666;
  wire[5:0] T935;
  wire[5:0] tgtPagesOH_44;
  wire[7:0] T936;
  wire[2:0] T937;
  wire[1:0] T938;
  wire T939;
  wire[7:0] T940;
  wire[7:0] T1667;
  wire[5:0] T941;
  wire[5:0] tgtPagesOH_45;
  wire[7:0] T942;
  wire[2:0] T943;
  wire T944;
  wire[7:0] T945;
  wire[7:0] T1668;
  wire[5:0] T946;
  wire[5:0] tgtPagesOH_46;
  wire[7:0] T947;
  wire[2:0] T948;
  wire[14:0] T949;
  wire[7:0] T950;
  wire[3:0] T951;
  wire[1:0] T952;
  wire T953;
  wire[7:0] T954;
  wire[7:0] T1669;
  wire[5:0] T955;
  wire[5:0] tgtPagesOH_47;
  wire[7:0] T956;
  wire[2:0] T957;
  wire T958;
  wire[7:0] T959;
  wire[7:0] T1670;
  wire[5:0] T960;
  wire[5:0] tgtPagesOH_48;
  wire[7:0] T961;
  wire[2:0] T962;
  wire[1:0] T963;
  wire T964;
  wire[7:0] T965;
  wire[7:0] T1671;
  wire[5:0] T966;
  wire[5:0] tgtPagesOH_49;
  wire[7:0] T967;
  wire[2:0] T968;
  wire T969;
  wire[7:0] T970;
  wire[7:0] T1672;
  wire[5:0] T971;
  wire[5:0] tgtPagesOH_50;
  wire[7:0] T972;
  wire[2:0] T973;
  wire[3:0] T974;
  wire[1:0] T975;
  wire T976;
  wire[7:0] T977;
  wire[7:0] T1673;
  wire[5:0] T978;
  wire[5:0] tgtPagesOH_51;
  wire[7:0] T979;
  wire[2:0] T980;
  wire T981;
  wire[7:0] T982;
  wire[7:0] T1674;
  wire[5:0] T983;
  wire[5:0] tgtPagesOH_52;
  wire[7:0] T984;
  wire[2:0] T985;
  wire[1:0] T986;
  wire T987;
  wire[7:0] T988;
  wire[7:0] T1675;
  wire[5:0] T989;
  wire[5:0] tgtPagesOH_53;
  wire[7:0] T990;
  wire[2:0] T991;
  wire T992;
  wire[7:0] T993;
  wire[7:0] T1676;
  wire[5:0] T994;
  wire[5:0] tgtPagesOH_54;
  wire[7:0] T995;
  wire[2:0] T996;
  wire[6:0] T997;
  wire[3:0] T998;
  wire[1:0] T999;
  wire T1000;
  wire[7:0] T1001;
  wire[7:0] T1677;
  wire[5:0] T1002;
  wire[5:0] tgtPagesOH_55;
  wire[7:0] T1003;
  wire[2:0] T1004;
  wire T1005;
  wire[7:0] T1006;
  wire[7:0] T1678;
  wire[5:0] T1007;
  wire[5:0] tgtPagesOH_56;
  wire[7:0] T1008;
  wire[2:0] T1009;
  wire[1:0] T1010;
  wire T1011;
  wire[7:0] T1012;
  wire[7:0] T1679;
  wire[5:0] T1013;
  wire[5:0] tgtPagesOH_57;
  wire[7:0] T1014;
  wire[2:0] T1015;
  wire T1016;
  wire[7:0] T1017;
  wire[7:0] T1680;
  wire[5:0] T1018;
  wire[5:0] tgtPagesOH_58;
  wire[7:0] T1019;
  wire[2:0] T1020;
  wire[2:0] T1021;
  wire[1:0] T1022;
  wire T1023;
  wire[7:0] T1024;
  wire[7:0] T1681;
  wire[5:0] T1025;
  wire[5:0] tgtPagesOH_59;
  wire[7:0] T1026;
  wire[2:0] T1027;
  wire T1028;
  wire[7:0] T1029;
  wire[7:0] T1682;
  wire[5:0] T1030;
  wire[5:0] tgtPagesOH_60;
  wire[7:0] T1031;
  wire[2:0] T1032;
  wire T1033;
  wire[7:0] T1034;
  wire[7:0] T1683;
  wire[5:0] T1035;
  wire[5:0] tgtPagesOH_61;
  wire[7:0] T1036;
  wire[2:0] T1037;
  wire[63:0] T1038;
  wire[63:0] T1039;
  wire[63:0] T1040;
  wire[63:0] T1684;
  wire[61:0] T1041;
  wire[63:0] T1042;
  wire[63:0] T1685;
  wire T1043;
  wire T1044;
  wire[63:0] T1045;
  wire[63:0] T1046;
  wire[63:0] T1686;
  wire T1047;
  wire T1048;
  wire[6:0] T1049;
  wire[5:0] T1050;
  wire T1051;
  wire[6:0] T1052;
  wire[6:0] T1053;
  wire[5:0] T1687;
  wire[4:0] T1688;
  wire[3:0] T1689;
  wire[2:0] T1690;
  wire[1:0] T1691;
  wire T1692;
  wire[1:0] T1693;
  wire[1:0] T1694;
  wire[3:0] T1695;
  wire[3:0] T1696;
  wire[7:0] T1697;
  wire[7:0] T1698;
  wire[15:0] T1699;
  wire[15:0] T1700;
  wire[31:0] T1701;
  wire[31:0] T1702;
  wire[29:0] T1703;
  wire[15:0] T1704;
  wire[7:0] T1705;
  wire[3:0] T1706;
  wire[1:0] T1707;
  wire T1708;
  wire T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[42:0] T1055;
  wire[42:0] T1056;
  wire[42:0] T1057;
  wire[12:0] T1058;
  wire[12:0] T1059;
  wire[12:0] T1060;
  reg [12:0] tgts [61:0];
  wire[12:0] T1061;
  wire[12:0] T1713;
  wire T1062;
  wire T1063;
  wire T1064;
  wire[12:0] T1065;
  wire[12:0] T1066;
  wire[12:0] T1067;
  wire T1068;
  wire[12:0] T1069;
  wire[12:0] T1070;
  wire[12:0] T1071;
  wire T1072;
  wire[12:0] T1073;
  wire[12:0] T1074;
  wire[12:0] T1075;
  wire T1076;
  wire[12:0] T1077;
  wire[12:0] T1078;
  wire[12:0] T1079;
  wire T1080;
  wire[12:0] T1081;
  wire[12:0] T1082;
  wire[12:0] T1083;
  wire T1084;
  wire[12:0] T1085;
  wire[12:0] T1086;
  wire[12:0] T1087;
  wire T1088;
  wire[12:0] T1089;
  wire[12:0] T1090;
  wire[12:0] T1091;
  wire T1092;
  wire[12:0] T1093;
  wire[12:0] T1094;
  wire[12:0] T1095;
  wire T1096;
  wire[12:0] T1097;
  wire[12:0] T1098;
  wire[12:0] T1099;
  wire T1100;
  wire[12:0] T1101;
  wire[12:0] T1102;
  wire[12:0] T1103;
  wire T1104;
  wire[12:0] T1105;
  wire[12:0] T1106;
  wire[12:0] T1107;
  wire T1108;
  wire[12:0] T1109;
  wire[12:0] T1110;
  wire[12:0] T1111;
  wire T1112;
  wire[12:0] T1113;
  wire[12:0] T1114;
  wire[12:0] T1115;
  wire T1116;
  wire[12:0] T1117;
  wire[12:0] T1118;
  wire[12:0] T1119;
  wire T1120;
  wire[12:0] T1121;
  wire[12:0] T1122;
  wire[12:0] T1123;
  wire T1124;
  wire[12:0] T1125;
  wire[12:0] T1126;
  wire[12:0] T1127;
  wire T1128;
  wire[12:0] T1129;
  wire[12:0] T1130;
  wire[12:0] T1131;
  wire T1132;
  wire[12:0] T1133;
  wire[12:0] T1134;
  wire[12:0] T1135;
  wire T1136;
  wire[12:0] T1137;
  wire[12:0] T1138;
  wire[12:0] T1139;
  wire T1140;
  wire[12:0] T1141;
  wire[12:0] T1142;
  wire[12:0] T1143;
  wire T1144;
  wire[12:0] T1145;
  wire[12:0] T1146;
  wire[12:0] T1147;
  wire T1148;
  wire[12:0] T1149;
  wire[12:0] T1150;
  wire[12:0] T1151;
  wire T1152;
  wire[12:0] T1153;
  wire[12:0] T1154;
  wire[12:0] T1155;
  wire T1156;
  wire[12:0] T1157;
  wire[12:0] T1158;
  wire[12:0] T1159;
  wire T1160;
  wire[12:0] T1161;
  wire[12:0] T1162;
  wire[12:0] T1163;
  wire T1164;
  wire[12:0] T1165;
  wire[12:0] T1166;
  wire[12:0] T1167;
  wire T1168;
  wire[12:0] T1169;
  wire[12:0] T1170;
  wire[12:0] T1171;
  wire T1172;
  wire[12:0] T1173;
  wire[12:0] T1174;
  wire[12:0] T1175;
  wire T1176;
  wire[12:0] T1177;
  wire[12:0] T1178;
  wire[12:0] T1179;
  wire T1180;
  wire[12:0] T1181;
  wire[12:0] T1182;
  wire[12:0] T1183;
  wire T1184;
  wire[12:0] T1185;
  wire[12:0] T1186;
  wire[12:0] T1187;
  wire T1188;
  wire[12:0] T1189;
  wire[12:0] T1190;
  wire[12:0] T1191;
  wire T1192;
  wire[12:0] T1193;
  wire[12:0] T1194;
  wire[12:0] T1195;
  wire T1196;
  wire[12:0] T1197;
  wire[12:0] T1198;
  wire[12:0] T1199;
  wire T1200;
  wire[12:0] T1201;
  wire[12:0] T1202;
  wire[12:0] T1203;
  wire T1204;
  wire[12:0] T1205;
  wire[12:0] T1206;
  wire[12:0] T1207;
  wire T1208;
  wire[12:0] T1209;
  wire[12:0] T1210;
  wire[12:0] T1211;
  wire T1212;
  wire[12:0] T1213;
  wire[12:0] T1214;
  wire[12:0] T1215;
  wire T1216;
  wire[12:0] T1217;
  wire[12:0] T1218;
  wire[12:0] T1219;
  wire T1220;
  wire[12:0] T1221;
  wire[12:0] T1222;
  wire[12:0] T1223;
  wire T1224;
  wire[12:0] T1225;
  wire[12:0] T1226;
  wire[12:0] T1227;
  wire T1228;
  wire[12:0] T1229;
  wire[12:0] T1230;
  wire[12:0] T1231;
  wire T1232;
  wire[12:0] T1233;
  wire[12:0] T1234;
  wire[12:0] T1235;
  wire T1236;
  wire[12:0] T1237;
  wire[12:0] T1238;
  wire[12:0] T1239;
  wire T1240;
  wire[12:0] T1241;
  wire[12:0] T1242;
  wire[12:0] T1243;
  wire T1244;
  wire[12:0] T1245;
  wire[12:0] T1246;
  wire[12:0] T1247;
  wire T1248;
  wire[12:0] T1249;
  wire[12:0] T1250;
  wire[12:0] T1251;
  wire T1252;
  wire[12:0] T1253;
  wire[12:0] T1254;
  wire[12:0] T1255;
  wire T1256;
  wire[12:0] T1257;
  wire[12:0] T1258;
  wire[12:0] T1259;
  wire T1260;
  wire[12:0] T1261;
  wire[12:0] T1262;
  wire[12:0] T1263;
  wire T1264;
  wire[12:0] T1265;
  wire[12:0] T1266;
  wire[12:0] T1267;
  wire T1268;
  wire[12:0] T1269;
  wire[12:0] T1270;
  wire[12:0] T1271;
  wire T1272;
  wire[12:0] T1273;
  wire[12:0] T1274;
  wire[12:0] T1275;
  wire T1276;
  wire[12:0] T1277;
  wire[12:0] T1278;
  wire[12:0] T1279;
  wire T1280;
  wire[12:0] T1281;
  wire[12:0] T1282;
  wire[12:0] T1283;
  wire T1284;
  wire[12:0] T1285;
  wire[12:0] T1286;
  wire[12:0] T1287;
  wire T1288;
  wire[12:0] T1289;
  wire[12:0] T1290;
  wire[12:0] T1291;
  wire T1292;
  wire[12:0] T1293;
  wire[12:0] T1294;
  wire[12:0] T1295;
  wire T1296;
  wire[12:0] T1297;
  wire[12:0] T1298;
  wire[12:0] T1299;
  wire T1300;
  wire[12:0] T1301;
  wire[12:0] T1302;
  wire[12:0] T1303;
  wire T1304;
  wire[12:0] T1305;
  wire[12:0] T1306;
  wire T1307;
  wire[29:0] T1308;
  wire[29:0] T1309;
  wire[29:0] T1310;
  wire T1311;
  wire[5:0] T1312;
  wire[5:0] T1313;
  wire T1314;
  wire[5:0] T1315;
  wire[5:0] T1316;
  wire T1317;
  wire[5:0] T1318;
  wire[5:0] T1319;
  wire T1320;
  wire[5:0] T1321;
  wire[5:0] T1322;
  wire T1323;
  wire[5:0] T1324;
  wire[5:0] T1325;
  wire T1326;
  wire[5:0] T1327;
  wire[5:0] T1328;
  wire T1329;
  wire[5:0] T1330;
  wire[5:0] T1331;
  wire T1332;
  wire[5:0] T1333;
  wire[5:0] T1334;
  wire T1335;
  wire[5:0] T1336;
  wire[5:0] T1337;
  wire T1338;
  wire[5:0] T1339;
  wire[5:0] T1340;
  wire T1341;
  wire[5:0] T1342;
  wire[5:0] T1343;
  wire T1344;
  wire[5:0] T1345;
  wire[5:0] T1346;
  wire T1347;
  wire[5:0] T1348;
  wire[5:0] T1349;
  wire T1350;
  wire[5:0] T1351;
  wire[5:0] T1352;
  wire T1353;
  wire[5:0] T1354;
  wire[5:0] T1355;
  wire T1356;
  wire[5:0] T1357;
  wire[5:0] T1358;
  wire T1359;
  wire[5:0] T1360;
  wire[5:0] T1361;
  wire T1362;
  wire[5:0] T1363;
  wire[5:0] T1364;
  wire T1365;
  wire[5:0] T1366;
  wire[5:0] T1367;
  wire T1368;
  wire[5:0] T1369;
  wire[5:0] T1370;
  wire T1371;
  wire[5:0] T1372;
  wire[5:0] T1373;
  wire T1374;
  wire[5:0] T1375;
  wire[5:0] T1376;
  wire T1377;
  wire[5:0] T1378;
  wire[5:0] T1379;
  wire T1380;
  wire[5:0] T1381;
  wire[5:0] T1382;
  wire T1383;
  wire[5:0] T1384;
  wire[5:0] T1385;
  wire T1386;
  wire[5:0] T1387;
  wire[5:0] T1388;
  wire T1389;
  wire[5:0] T1390;
  wire[5:0] T1391;
  wire T1392;
  wire[5:0] T1393;
  wire[5:0] T1394;
  wire T1395;
  wire[5:0] T1396;
  wire[5:0] T1397;
  wire T1398;
  wire[5:0] T1399;
  wire[5:0] T1400;
  wire T1401;
  wire[5:0] T1402;
  wire[5:0] T1403;
  wire T1404;
  wire[5:0] T1405;
  wire[5:0] T1406;
  wire T1407;
  wire[5:0] T1408;
  wire[5:0] T1409;
  wire T1410;
  wire[5:0] T1411;
  wire[5:0] T1412;
  wire T1413;
  wire[5:0] T1414;
  wire[5:0] T1415;
  wire T1416;
  wire[5:0] T1417;
  wire[5:0] T1418;
  wire T1419;
  wire[5:0] T1420;
  wire[5:0] T1421;
  wire T1422;
  wire[5:0] T1423;
  wire[5:0] T1424;
  wire T1425;
  wire[5:0] T1426;
  wire[5:0] T1427;
  wire T1428;
  wire[5:0] T1429;
  wire[5:0] T1430;
  wire T1431;
  wire[5:0] T1432;
  wire[5:0] T1433;
  wire T1434;
  wire[5:0] T1435;
  wire[5:0] T1436;
  wire T1437;
  wire[5:0] T1438;
  wire[5:0] T1439;
  wire T1440;
  wire[5:0] T1441;
  wire[5:0] T1442;
  wire T1443;
  wire[5:0] T1444;
  wire[5:0] T1445;
  wire T1446;
  wire[5:0] T1447;
  wire[5:0] T1448;
  wire T1449;
  wire[5:0] T1450;
  wire[5:0] T1451;
  wire T1452;
  wire[5:0] T1453;
  wire[5:0] T1454;
  wire T1455;
  wire[5:0] T1456;
  wire[5:0] T1457;
  wire T1458;
  wire[5:0] T1459;
  wire[5:0] T1460;
  wire T1461;
  wire[5:0] T1462;
  wire[5:0] T1463;
  wire T1464;
  wire[5:0] T1465;
  wire[5:0] T1466;
  wire T1467;
  wire[5:0] T1468;
  wire[5:0] T1469;
  wire T1470;
  wire[5:0] T1471;
  wire[5:0] T1472;
  wire T1473;
  wire[5:0] T1474;
  wire[5:0] T1475;
  wire T1476;
  wire[5:0] T1477;
  wire[5:0] T1478;
  wire T1479;
  wire[5:0] T1480;
  wire[5:0] T1481;
  wire T1482;
  wire[5:0] T1483;
  wire[5:0] T1484;
  wire T1485;
  wire[5:0] T1486;
  wire[5:0] T1487;
  wire T1488;
  wire[5:0] T1489;
  wire[5:0] T1490;
  wire T1491;
  wire[5:0] T1492;
  wire[5:0] T1493;
  wire T1494;
  wire[5:0] T1495;
  wire T1496;
  wire[29:0] T1497;
  wire[29:0] T1498;
  wire[29:0] T1499;
  wire T1500;
  wire[29:0] T1501;
  wire[29:0] T1502;
  wire[29:0] T1503;
  wire T1504;
  wire[29:0] T1505;
  wire[29:0] T1506;
  wire[29:0] T1507;
  wire T1508;
  wire[29:0] T1509;
  wire[29:0] T1510;
  wire[29:0] T1511;
  wire T1512;
  wire[29:0] T1513;
  wire[29:0] T1514;
  wire T1515;
  wire[42:0] T1516;
  reg [42:0] R1517;
  wire[42:0] T1518;
  wire T1519;
  wire T1520;
  wire[1:0] T1521;
  wire T1522;
  wire T1523;
  reg  R1524;
  wire T1714;
  wire T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  reg [1:0] R1531;
  wire[1:0] T1715;
  wire[1:0] T1532;
  wire[1:0] T1533;
  wire[1:0] T1534;
  wire[1:0] T1535;
  wire T1536;
  wire T1537;
  wire[1:0] T1538;
  wire T1539;
  wire T1540;
  wire T1541;
  wire T1542;
  wire T1543;
  reg [42:0] R1544;
  wire[42:0] T1545;
  wire T1546;
  wire T1547;
  wire T1548;
  wire T1549;
  wire T1550;
  wire[61:0] T1551;
  reg [61:0] useRAS;
  wire[61:0] T1716;
  wire[63:0] T1552;
  wire[63:0] T1717;
  wire[63:0] T1553;
  wire[63:0] T1554;
  wire[63:0] T1555;
  wire[63:0] T1718;
  wire[61:0] T1556;
  wire[63:0] T1557;
  wire[63:0] T1719;
  wire T1558;
  wire T1559;
  reg  R1560;
  wire T1561;
  wire[63:0] T1562;
  wire[63:0] T1563;
  wire[63:0] T1720;
  wire T1564;
  wire T1565;
  wire T1566;
  wire T1567;
  reg [0:0] brIdx [61:0];
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire[61:0] T1575;
  wire T1576;
  wire T1577;
  wire T1578;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R7 = {1{$random}};
    for (initvar = 0; initvar < 128; initvar = initvar+1)
      T10[initvar] = {1{$random}};
    R25 = {1{$random}};
    isJump = {2{$random}};
    R42 = {1{$random}};
    R49 = {1{$random}};
    updateHit = {1{$random}};
    R54 = {1{$random}};
    pageValid = {1{$random}};
    R75 = {1{$random}};
    R87 = {2{$random}};
    for (initvar = 0; initvar < 6; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {2{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R1517 = {2{$random}};
    R1524 = {1{$random}};
    R1531 = {1{$random}};
    R1544 = {2{$random}};
    useRAS = {2{$random}};
    R1560 = {1{$random}};
    for (initvar = 0; initvar < 62; initvar = initvar+1)
      brIdx[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_btb_update_valid ? io_btb_update_bits_target : R4;
  assign T6 = R7 ^ 1'h1;
  assign T1579 = reset ? 1'h0 : io_btb_update_valid;
  assign io_resp_bits_bht_value = T8;
  assign T8 = T9;
  assign T9 = T10[T24];
  assign T12 = {io_bht_update_bits_taken, T13};
  assign T13 = T18 | T14;
  assign T14 = T15 & io_bht_update_bits_taken;
  assign T15 = T17 | T16;
  assign T16 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T17 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T18 = T20 & T19;
  assign T19 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T20 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T21 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T22 = T23 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T23 = io_bht_update_bits_pc[4'h8:2'h2];
  assign T24 = T1052 ^ R25;
  assign T26 = T1051 ? T1049 : T27;
  assign T27 = T31 ? T28 : R25;
  assign T28 = {T30, T29};
  assign T29 = R25[3'h6:1'h1];
  assign T30 = T8[1'h0:1'h0];
  assign T31 = T1047 & T32;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T34 != 62'h0;
  assign T34 = hits & isJump;
  assign T1580 = T35[6'h3d:1'h0];
  assign T35 = R7 ? T36 : T1581;
  assign T1581 = {2'h0, isJump};
  assign T36 = T56 | T37;
  assign T37 = T1584 & T38;
  assign T38 = T40 | T1582;
  assign T1582 = {2'h0, T39};
  assign T39 = isJump ^ isJump;
  assign T40 = 1'h1 << T41;
  assign T41 = updateHit ? R49 : R42;
  assign T1583 = reset ? 6'h0 : T43;
  assign T43 = T47 ? T44 : R42;
  assign T44 = T46 ? 6'h0 : T45;
  assign T45 = R42 + 6'h1;
  assign T46 = R42 == 6'h3d;
  assign T47 = R7 & T48;
  assign T48 = updateHit ^ 1'h1;
  assign T50 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : R49;
  assign T51 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : updateHit;
  assign T1584 = T52 ? 64'hffffffffffffffff : 64'h0;
  assign T52 = T53;
  assign T53 = R54;
  assign T55 = io_btb_update_valid ? io_btb_update_bits_isJump : R54;
  assign T56 = T1585 & T57;
  assign T57 = ~ T38;
  assign T1585 = {2'h0, isJump};
  assign hits = T466 & T58;
  assign T58 = T59;
  assign T59 = {T312, T60};
  assign T60 = {T238, T61};
  assign T61 = {T199, T62};
  assign T62 = {T180, T63};
  assign T63 = {T171, T64};
  assign T64 = {T167, T65};
  assign T65 = T66 != 6'h0;
  assign T66 = idxPagesOH_0 & pageHit;
  assign pageHit = T143 & pageValid;
  assign T1586 = T1587[3'h5:1'h0];
  assign T1587 = reset ? 8'h0 : T67;
  assign T67 = io_invalidate ? 8'h0 : T68;
  assign T68 = T142 ? T69 : T1588;
  assign T1588 = {2'h0, pageValid};
  assign T69 = T1594 | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T1589;
  assign T1589 = {2'h0, T70};
  assign T70 = T72 | T1590;
  assign T1590 = {5'h0, T71};
  assign T71 = idxPageUpdateOH[3'h5:3'h5];
  assign T72 = T73 << 1'h1;
  assign T73 = idxPageUpdateOH[3'h4:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? T1592 : idxPageRepl;
  assign idxPageRepl = T74;
  assign T74 = 1'h1 << R75;
  assign T1591 = reset ? 3'h0 : T76;
  assign T76 = T80 ? T77 : R75;
  assign T77 = T79 ? 3'h0 : T78;
  assign T78 = R75 + 3'h1;
  assign T79 = R75 == 3'h5;
  assign T80 = R7 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = useUpdatePageHit ^ 1'h1;
  assign T1592 = {2'h0, updatePageHit};
  assign updatePageHit = T81 & pageValid;
  assign T81 = T82;
  assign T82 = {T128, T83};
  assign T83 = {T126, T84};
  assign T84 = {T124, T85};
  assign T85 = T89 == T86;
  assign T86 = R87 >> 4'hd;
  assign T88 = io_btb_update_valid ? io_btb_update_bits_pc : R87;
  assign T89 = pages[3'h0];
  assign T91 = T94 ? T93 : T92;
  assign T92 = R87 >> 4'hd;
  assign T93 = io_req_bits_addr >> 4'hd;
  assign T94 = T95 != 8'h0;
  assign T95 = idxPageUpdateOH & 8'h15;
  assign T96 = R7 & T97;
  assign T97 = T99 & T98;
  assign T98 = pageReplEn[3'h5:3'h5];
  assign T99 = T94 ? doTgtPageRepl : doIdxPageRepl;
  assign T101 = R7 & T102;
  assign T102 = T99 & T103;
  assign T103 = pageReplEn[2'h3:2'h3];
  assign T105 = R7 & T106;
  assign T106 = T99 & T107;
  assign T107 = pageReplEn[1'h1:1'h1];
  assign T109 = T94 ? T111 : T110;
  assign T110 = io_req_bits_addr >> 4'hd;
  assign T111 = R87 >> 4'hd;
  assign T112 = R7 & T113;
  assign T113 = T115 & T114;
  assign T114 = pageReplEn[3'h4:3'h4];
  assign T115 = T94 ? doIdxPageRepl : doTgtPageRepl;
  assign T117 = R7 & T118;
  assign T118 = T115 & T119;
  assign T119 = pageReplEn[2'h2:2'h2];
  assign T121 = R7 & T122;
  assign T122 = T115 & T123;
  assign T123 = pageReplEn[1'h0:1'h0];
  assign T124 = T125 == T86;
  assign T125 = pages[3'h1];
  assign T126 = T127 == T86;
  assign T127 = pages[3'h2];
  assign T128 = {T134, T129};
  assign T129 = {T132, T130};
  assign T130 = T131 == T86;
  assign T131 = pages[3'h3];
  assign T132 = T133 == T86;
  assign T133 = pages[3'h4];
  assign T134 = T135 == T86;
  assign T135 = pages[3'h5];
  assign useUpdatePageHit = updatePageHit != 6'h0;
  assign samePage = T137 == T136;
  assign T136 = io_req_bits_addr >> 4'hd;
  assign T137 = R87 >> 4'hd;
  assign doTgtPageRepl = T141 & T138;
  assign T138 = usePageHit ^ 1'h1;
  assign usePageHit = T139 != 8'h0;
  assign T139 = T1593 & T140;
  assign T140 = ~ idxPageReplEn;
  assign T1593 = {2'h0, pageHit};
  assign T141 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0;
  assign T1594 = {2'h0, pageValid};
  assign T142 = R7 & doPageRepl;
  assign T143 = T144;
  assign T144 = {T154, T145};
  assign T145 = {T152, T146};
  assign T146 = {T150, T147};
  assign T147 = T149 == T148;
  assign T148 = io_req_bits_addr >> 4'hd;
  assign T149 = pages[3'h0];
  assign T150 = T151 == T148;
  assign T151 = pages[3'h1];
  assign T152 = T153 == T148;
  assign T153 = pages[3'h2];
  assign T154 = {T160, T155};
  assign T155 = {T158, T156};
  assign T156 = T157 == T148;
  assign T157 = pages[3'h3];
  assign T158 = T159 == T148;
  assign T159 = pages[3'h4];
  assign T160 = T161 == T148;
  assign T161 = pages[3'h5];
  assign idxPagesOH_0 = T162[3'h5:1'h0];
  assign T162 = 1'h1 << T163;
  assign T163 = idxPages[6'h0];
  assign T1595 = {T1605, T1596};
  assign T1596 = {T1604, T1597};
  assign T1597 = T1598[1'h1:1'h1];
  assign T1598 = T1603 | T1599;
  assign T1599 = T1600[1'h1:1'h0];
  assign T1600 = T1602 | T1601;
  assign T1601 = idxPageUpdateOH[2'h3:1'h0];
  assign T1602 = idxPageUpdateOH[3'h7:3'h4];
  assign T1603 = T1600[2'h3:2'h2];
  assign T1604 = T1603 != 2'h0;
  assign T1605 = T1602 != 4'h0;
  assign T165 = R7 & T166;
  assign T166 = T41 < 6'h3e;
  assign T167 = T168 != 6'h0;
  assign T168 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T169[3'h5:1'h0];
  assign T169 = 1'h1 << T170;
  assign T170 = idxPages[6'h1];
  assign T171 = {T176, T172};
  assign T172 = T173 != 6'h0;
  assign T173 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T174[3'h5:1'h0];
  assign T174 = 1'h1 << T175;
  assign T175 = idxPages[6'h2];
  assign T176 = T177 != 6'h0;
  assign T177 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T178[3'h5:1'h0];
  assign T178 = 1'h1 << T179;
  assign T179 = idxPages[6'h3];
  assign T180 = {T190, T181};
  assign T181 = {T186, T182};
  assign T182 = T183 != 6'h0;
  assign T183 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T184[3'h5:1'h0];
  assign T184 = 1'h1 << T185;
  assign T185 = idxPages[6'h4];
  assign T186 = T187 != 6'h0;
  assign T187 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T188[3'h5:1'h0];
  assign T188 = 1'h1 << T189;
  assign T189 = idxPages[6'h5];
  assign T190 = {T195, T191};
  assign T191 = T192 != 6'h0;
  assign T192 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T193[3'h5:1'h0];
  assign T193 = 1'h1 << T194;
  assign T194 = idxPages[6'h6];
  assign T195 = T196 != 6'h0;
  assign T196 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T197[3'h5:1'h0];
  assign T197 = 1'h1 << T198;
  assign T198 = idxPages[6'h7];
  assign T199 = {T219, T200};
  assign T200 = {T210, T201};
  assign T201 = {T206, T202};
  assign T202 = T203 != 6'h0;
  assign T203 = idxPagesOH_8 & pageHit;
  assign idxPagesOH_8 = T204[3'h5:1'h0];
  assign T204 = 1'h1 << T205;
  assign T205 = idxPages[6'h8];
  assign T206 = T207 != 6'h0;
  assign T207 = idxPagesOH_9 & pageHit;
  assign idxPagesOH_9 = T208[3'h5:1'h0];
  assign T208 = 1'h1 << T209;
  assign T209 = idxPages[6'h9];
  assign T210 = {T215, T211};
  assign T211 = T212 != 6'h0;
  assign T212 = idxPagesOH_10 & pageHit;
  assign idxPagesOH_10 = T213[3'h5:1'h0];
  assign T213 = 1'h1 << T214;
  assign T214 = idxPages[6'ha];
  assign T215 = T216 != 6'h0;
  assign T216 = idxPagesOH_11 & pageHit;
  assign idxPagesOH_11 = T217[3'h5:1'h0];
  assign T217 = 1'h1 << T218;
  assign T218 = idxPages[6'hb];
  assign T219 = {T229, T220};
  assign T220 = {T225, T221};
  assign T221 = T222 != 6'h0;
  assign T222 = idxPagesOH_12 & pageHit;
  assign idxPagesOH_12 = T223[3'h5:1'h0];
  assign T223 = 1'h1 << T224;
  assign T224 = idxPages[6'hc];
  assign T225 = T226 != 6'h0;
  assign T226 = idxPagesOH_13 & pageHit;
  assign idxPagesOH_13 = T227[3'h5:1'h0];
  assign T227 = 1'h1 << T228;
  assign T228 = idxPages[6'hd];
  assign T229 = {T234, T230};
  assign T230 = T231 != 6'h0;
  assign T231 = idxPagesOH_14 & pageHit;
  assign idxPagesOH_14 = T232[3'h5:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = idxPages[6'he];
  assign T234 = T235 != 6'h0;
  assign T235 = idxPagesOH_15 & pageHit;
  assign idxPagesOH_15 = T236[3'h5:1'h0];
  assign T236 = 1'h1 << T237;
  assign T237 = idxPages[6'hf];
  assign T238 = {T278, T239};
  assign T239 = {T259, T240};
  assign T240 = {T250, T241};
  assign T241 = {T246, T242};
  assign T242 = T243 != 6'h0;
  assign T243 = idxPagesOH_16 & pageHit;
  assign idxPagesOH_16 = T244[3'h5:1'h0];
  assign T244 = 1'h1 << T245;
  assign T245 = idxPages[6'h10];
  assign T246 = T247 != 6'h0;
  assign T247 = idxPagesOH_17 & pageHit;
  assign idxPagesOH_17 = T248[3'h5:1'h0];
  assign T248 = 1'h1 << T249;
  assign T249 = idxPages[6'h11];
  assign T250 = {T255, T251};
  assign T251 = T252 != 6'h0;
  assign T252 = idxPagesOH_18 & pageHit;
  assign idxPagesOH_18 = T253[3'h5:1'h0];
  assign T253 = 1'h1 << T254;
  assign T254 = idxPages[6'h12];
  assign T255 = T256 != 6'h0;
  assign T256 = idxPagesOH_19 & pageHit;
  assign idxPagesOH_19 = T257[3'h5:1'h0];
  assign T257 = 1'h1 << T258;
  assign T258 = idxPages[6'h13];
  assign T259 = {T269, T260};
  assign T260 = {T265, T261};
  assign T261 = T262 != 6'h0;
  assign T262 = idxPagesOH_20 & pageHit;
  assign idxPagesOH_20 = T263[3'h5:1'h0];
  assign T263 = 1'h1 << T264;
  assign T264 = idxPages[6'h14];
  assign T265 = T266 != 6'h0;
  assign T266 = idxPagesOH_21 & pageHit;
  assign idxPagesOH_21 = T267[3'h5:1'h0];
  assign T267 = 1'h1 << T268;
  assign T268 = idxPages[6'h15];
  assign T269 = {T274, T270};
  assign T270 = T271 != 6'h0;
  assign T271 = idxPagesOH_22 & pageHit;
  assign idxPagesOH_22 = T272[3'h5:1'h0];
  assign T272 = 1'h1 << T273;
  assign T273 = idxPages[6'h16];
  assign T274 = T275 != 6'h0;
  assign T275 = idxPagesOH_23 & pageHit;
  assign idxPagesOH_23 = T276[3'h5:1'h0];
  assign T276 = 1'h1 << T277;
  assign T277 = idxPages[6'h17];
  assign T278 = {T298, T279};
  assign T279 = {T289, T280};
  assign T280 = {T285, T281};
  assign T281 = T282 != 6'h0;
  assign T282 = idxPagesOH_24 & pageHit;
  assign idxPagesOH_24 = T283[3'h5:1'h0];
  assign T283 = 1'h1 << T284;
  assign T284 = idxPages[6'h18];
  assign T285 = T286 != 6'h0;
  assign T286 = idxPagesOH_25 & pageHit;
  assign idxPagesOH_25 = T287[3'h5:1'h0];
  assign T287 = 1'h1 << T288;
  assign T288 = idxPages[6'h19];
  assign T289 = {T294, T290};
  assign T290 = T291 != 6'h0;
  assign T291 = idxPagesOH_26 & pageHit;
  assign idxPagesOH_26 = T292[3'h5:1'h0];
  assign T292 = 1'h1 << T293;
  assign T293 = idxPages[6'h1a];
  assign T294 = T295 != 6'h0;
  assign T295 = idxPagesOH_27 & pageHit;
  assign idxPagesOH_27 = T296[3'h5:1'h0];
  assign T296 = 1'h1 << T297;
  assign T297 = idxPages[6'h1b];
  assign T298 = {T308, T299};
  assign T299 = {T304, T300};
  assign T300 = T301 != 6'h0;
  assign T301 = idxPagesOH_28 & pageHit;
  assign idxPagesOH_28 = T302[3'h5:1'h0];
  assign T302 = 1'h1 << T303;
  assign T303 = idxPages[6'h1c];
  assign T304 = T305 != 6'h0;
  assign T305 = idxPagesOH_29 & pageHit;
  assign idxPagesOH_29 = T306[3'h5:1'h0];
  assign T306 = 1'h1 << T307;
  assign T307 = idxPages[6'h1d];
  assign T308 = T309 != 6'h0;
  assign T309 = idxPagesOH_30 & pageHit;
  assign idxPagesOH_30 = T310[3'h5:1'h0];
  assign T310 = 1'h1 << T311;
  assign T311 = idxPages[6'h1e];
  assign T312 = {T392, T313};
  assign T313 = {T353, T314};
  assign T314 = {T334, T315};
  assign T315 = {T325, T316};
  assign T316 = {T321, T317};
  assign T317 = T318 != 6'h0;
  assign T318 = idxPagesOH_31 & pageHit;
  assign idxPagesOH_31 = T319[3'h5:1'h0];
  assign T319 = 1'h1 << T320;
  assign T320 = idxPages[6'h1f];
  assign T321 = T322 != 6'h0;
  assign T322 = idxPagesOH_32 & pageHit;
  assign idxPagesOH_32 = T323[3'h5:1'h0];
  assign T323 = 1'h1 << T324;
  assign T324 = idxPages[6'h20];
  assign T325 = {T330, T326};
  assign T326 = T327 != 6'h0;
  assign T327 = idxPagesOH_33 & pageHit;
  assign idxPagesOH_33 = T328[3'h5:1'h0];
  assign T328 = 1'h1 << T329;
  assign T329 = idxPages[6'h21];
  assign T330 = T331 != 6'h0;
  assign T331 = idxPagesOH_34 & pageHit;
  assign idxPagesOH_34 = T332[3'h5:1'h0];
  assign T332 = 1'h1 << T333;
  assign T333 = idxPages[6'h22];
  assign T334 = {T344, T335};
  assign T335 = {T340, T336};
  assign T336 = T337 != 6'h0;
  assign T337 = idxPagesOH_35 & pageHit;
  assign idxPagesOH_35 = T338[3'h5:1'h0];
  assign T338 = 1'h1 << T339;
  assign T339 = idxPages[6'h23];
  assign T340 = T341 != 6'h0;
  assign T341 = idxPagesOH_36 & pageHit;
  assign idxPagesOH_36 = T342[3'h5:1'h0];
  assign T342 = 1'h1 << T343;
  assign T343 = idxPages[6'h24];
  assign T344 = {T349, T345};
  assign T345 = T346 != 6'h0;
  assign T346 = idxPagesOH_37 & pageHit;
  assign idxPagesOH_37 = T347[3'h5:1'h0];
  assign T347 = 1'h1 << T348;
  assign T348 = idxPages[6'h25];
  assign T349 = T350 != 6'h0;
  assign T350 = idxPagesOH_38 & pageHit;
  assign idxPagesOH_38 = T351[3'h5:1'h0];
  assign T351 = 1'h1 << T352;
  assign T352 = idxPages[6'h26];
  assign T353 = {T373, T354};
  assign T354 = {T364, T355};
  assign T355 = {T360, T356};
  assign T356 = T357 != 6'h0;
  assign T357 = idxPagesOH_39 & pageHit;
  assign idxPagesOH_39 = T358[3'h5:1'h0];
  assign T358 = 1'h1 << T359;
  assign T359 = idxPages[6'h27];
  assign T360 = T361 != 6'h0;
  assign T361 = idxPagesOH_40 & pageHit;
  assign idxPagesOH_40 = T362[3'h5:1'h0];
  assign T362 = 1'h1 << T363;
  assign T363 = idxPages[6'h28];
  assign T364 = {T369, T365};
  assign T365 = T366 != 6'h0;
  assign T366 = idxPagesOH_41 & pageHit;
  assign idxPagesOH_41 = T367[3'h5:1'h0];
  assign T367 = 1'h1 << T368;
  assign T368 = idxPages[6'h29];
  assign T369 = T370 != 6'h0;
  assign T370 = idxPagesOH_42 & pageHit;
  assign idxPagesOH_42 = T371[3'h5:1'h0];
  assign T371 = 1'h1 << T372;
  assign T372 = idxPages[6'h2a];
  assign T373 = {T383, T374};
  assign T374 = {T379, T375};
  assign T375 = T376 != 6'h0;
  assign T376 = idxPagesOH_43 & pageHit;
  assign idxPagesOH_43 = T377[3'h5:1'h0];
  assign T377 = 1'h1 << T378;
  assign T378 = idxPages[6'h2b];
  assign T379 = T380 != 6'h0;
  assign T380 = idxPagesOH_44 & pageHit;
  assign idxPagesOH_44 = T381[3'h5:1'h0];
  assign T381 = 1'h1 << T382;
  assign T382 = idxPages[6'h2c];
  assign T383 = {T388, T384};
  assign T384 = T385 != 6'h0;
  assign T385 = idxPagesOH_45 & pageHit;
  assign idxPagesOH_45 = T386[3'h5:1'h0];
  assign T386 = 1'h1 << T387;
  assign T387 = idxPages[6'h2d];
  assign T388 = T389 != 6'h0;
  assign T389 = idxPagesOH_46 & pageHit;
  assign idxPagesOH_46 = T390[3'h5:1'h0];
  assign T390 = 1'h1 << T391;
  assign T391 = idxPages[6'h2e];
  assign T392 = {T432, T393};
  assign T393 = {T413, T394};
  assign T394 = {T404, T395};
  assign T395 = {T400, T396};
  assign T396 = T397 != 6'h0;
  assign T397 = idxPagesOH_47 & pageHit;
  assign idxPagesOH_47 = T398[3'h5:1'h0];
  assign T398 = 1'h1 << T399;
  assign T399 = idxPages[6'h2f];
  assign T400 = T401 != 6'h0;
  assign T401 = idxPagesOH_48 & pageHit;
  assign idxPagesOH_48 = T402[3'h5:1'h0];
  assign T402 = 1'h1 << T403;
  assign T403 = idxPages[6'h30];
  assign T404 = {T409, T405};
  assign T405 = T406 != 6'h0;
  assign T406 = idxPagesOH_49 & pageHit;
  assign idxPagesOH_49 = T407[3'h5:1'h0];
  assign T407 = 1'h1 << T408;
  assign T408 = idxPages[6'h31];
  assign T409 = T410 != 6'h0;
  assign T410 = idxPagesOH_50 & pageHit;
  assign idxPagesOH_50 = T411[3'h5:1'h0];
  assign T411 = 1'h1 << T412;
  assign T412 = idxPages[6'h32];
  assign T413 = {T423, T414};
  assign T414 = {T419, T415};
  assign T415 = T416 != 6'h0;
  assign T416 = idxPagesOH_51 & pageHit;
  assign idxPagesOH_51 = T417[3'h5:1'h0];
  assign T417 = 1'h1 << T418;
  assign T418 = idxPages[6'h33];
  assign T419 = T420 != 6'h0;
  assign T420 = idxPagesOH_52 & pageHit;
  assign idxPagesOH_52 = T421[3'h5:1'h0];
  assign T421 = 1'h1 << T422;
  assign T422 = idxPages[6'h34];
  assign T423 = {T428, T424};
  assign T424 = T425 != 6'h0;
  assign T425 = idxPagesOH_53 & pageHit;
  assign idxPagesOH_53 = T426[3'h5:1'h0];
  assign T426 = 1'h1 << T427;
  assign T427 = idxPages[6'h35];
  assign T428 = T429 != 6'h0;
  assign T429 = idxPagesOH_54 & pageHit;
  assign idxPagesOH_54 = T430[3'h5:1'h0];
  assign T430 = 1'h1 << T431;
  assign T431 = idxPages[6'h36];
  assign T432 = {T452, T433};
  assign T433 = {T443, T434};
  assign T434 = {T439, T435};
  assign T435 = T436 != 6'h0;
  assign T436 = idxPagesOH_55 & pageHit;
  assign idxPagesOH_55 = T437[3'h5:1'h0];
  assign T437 = 1'h1 << T438;
  assign T438 = idxPages[6'h37];
  assign T439 = T440 != 6'h0;
  assign T440 = idxPagesOH_56 & pageHit;
  assign idxPagesOH_56 = T441[3'h5:1'h0];
  assign T441 = 1'h1 << T442;
  assign T442 = idxPages[6'h38];
  assign T443 = {T448, T444};
  assign T444 = T445 != 6'h0;
  assign T445 = idxPagesOH_57 & pageHit;
  assign idxPagesOH_57 = T446[3'h5:1'h0];
  assign T446 = 1'h1 << T447;
  assign T447 = idxPages[6'h39];
  assign T448 = T449 != 6'h0;
  assign T449 = idxPagesOH_58 & pageHit;
  assign idxPagesOH_58 = T450[3'h5:1'h0];
  assign T450 = 1'h1 << T451;
  assign T451 = idxPages[6'h3a];
  assign T452 = {T462, T453};
  assign T453 = {T458, T454};
  assign T454 = T455 != 6'h0;
  assign T455 = idxPagesOH_59 & pageHit;
  assign idxPagesOH_59 = T456[3'h5:1'h0];
  assign T456 = 1'h1 << T457;
  assign T457 = idxPages[6'h3b];
  assign T458 = T459 != 6'h0;
  assign T459 = idxPagesOH_60 & pageHit;
  assign idxPagesOH_60 = T460[3'h5:1'h0];
  assign T460 = 1'h1 << T461;
  assign T461 = idxPages[6'h3c];
  assign T462 = T463 != 6'h0;
  assign T463 = idxPagesOH_61 & pageHit;
  assign idxPagesOH_61 = T464[3'h5:1'h0];
  assign T464 = 1'h1 << T465;
  assign T465 = idxPages[6'h3d];
  assign T466 = idxValid & T467;
  assign T467 = T468;
  assign T468 = {T565, T469};
  assign T469 = {T521, T470};
  assign T470 = {T498, T471};
  assign T471 = {T487, T472};
  assign T472 = {T482, T473};
  assign T473 = {T480, T474};
  assign T474 = T476 == T475;
  assign T475 = io_req_bits_addr[4'hc:1'h0];
  assign T476 = idxs[6'h0];
  assign T1606 = R87[4'hc:1'h0];
  assign T478 = R7 & T479;
  assign T479 = T41 < 6'h3e;
  assign T480 = T481 == T475;
  assign T481 = idxs[6'h1];
  assign T482 = {T485, T483};
  assign T483 = T484 == T475;
  assign T484 = idxs[6'h2];
  assign T485 = T486 == T475;
  assign T486 = idxs[6'h3];
  assign T487 = {T493, T488};
  assign T488 = {T491, T489};
  assign T489 = T490 == T475;
  assign T490 = idxs[6'h4];
  assign T491 = T492 == T475;
  assign T492 = idxs[6'h5];
  assign T493 = {T496, T494};
  assign T494 = T495 == T475;
  assign T495 = idxs[6'h6];
  assign T496 = T497 == T475;
  assign T497 = idxs[6'h7];
  assign T498 = {T510, T499};
  assign T499 = {T505, T500};
  assign T500 = {T503, T501};
  assign T501 = T502 == T475;
  assign T502 = idxs[6'h8];
  assign T503 = T504 == T475;
  assign T504 = idxs[6'h9];
  assign T505 = {T508, T506};
  assign T506 = T507 == T475;
  assign T507 = idxs[6'ha];
  assign T508 = T509 == T475;
  assign T509 = idxs[6'hb];
  assign T510 = {T516, T511};
  assign T511 = {T514, T512};
  assign T512 = T513 == T475;
  assign T513 = idxs[6'hc];
  assign T514 = T515 == T475;
  assign T515 = idxs[6'hd];
  assign T516 = {T519, T517};
  assign T517 = T518 == T475;
  assign T518 = idxs[6'he];
  assign T519 = T520 == T475;
  assign T520 = idxs[6'hf];
  assign T521 = {T545, T522};
  assign T522 = {T534, T523};
  assign T523 = {T529, T524};
  assign T524 = {T527, T525};
  assign T525 = T526 == T475;
  assign T526 = idxs[6'h10];
  assign T527 = T528 == T475;
  assign T528 = idxs[6'h11];
  assign T529 = {T532, T530};
  assign T530 = T531 == T475;
  assign T531 = idxs[6'h12];
  assign T532 = T533 == T475;
  assign T533 = idxs[6'h13];
  assign T534 = {T540, T535};
  assign T535 = {T538, T536};
  assign T536 = T537 == T475;
  assign T537 = idxs[6'h14];
  assign T538 = T539 == T475;
  assign T539 = idxs[6'h15];
  assign T540 = {T543, T541};
  assign T541 = T542 == T475;
  assign T542 = idxs[6'h16];
  assign T543 = T544 == T475;
  assign T544 = idxs[6'h17];
  assign T545 = {T557, T546};
  assign T546 = {T552, T547};
  assign T547 = {T550, T548};
  assign T548 = T549 == T475;
  assign T549 = idxs[6'h18];
  assign T550 = T551 == T475;
  assign T551 = idxs[6'h19];
  assign T552 = {T555, T553};
  assign T553 = T554 == T475;
  assign T554 = idxs[6'h1a];
  assign T555 = T556 == T475;
  assign T556 = idxs[6'h1b];
  assign T557 = {T563, T558};
  assign T558 = {T561, T559};
  assign T559 = T560 == T475;
  assign T560 = idxs[6'h1c];
  assign T561 = T562 == T475;
  assign T562 = idxs[6'h1d];
  assign T563 = T564 == T475;
  assign T564 = idxs[6'h1e];
  assign T565 = {T613, T566};
  assign T566 = {T590, T567};
  assign T567 = {T579, T568};
  assign T568 = {T574, T569};
  assign T569 = {T572, T570};
  assign T570 = T571 == T475;
  assign T571 = idxs[6'h1f];
  assign T572 = T573 == T475;
  assign T573 = idxs[6'h20];
  assign T574 = {T577, T575};
  assign T575 = T576 == T475;
  assign T576 = idxs[6'h21];
  assign T577 = T578 == T475;
  assign T578 = idxs[6'h22];
  assign T579 = {T585, T580};
  assign T580 = {T583, T581};
  assign T581 = T582 == T475;
  assign T582 = idxs[6'h23];
  assign T583 = T584 == T475;
  assign T584 = idxs[6'h24];
  assign T585 = {T588, T586};
  assign T586 = T587 == T475;
  assign T587 = idxs[6'h25];
  assign T588 = T589 == T475;
  assign T589 = idxs[6'h26];
  assign T590 = {T602, T591};
  assign T591 = {T597, T592};
  assign T592 = {T595, T593};
  assign T593 = T594 == T475;
  assign T594 = idxs[6'h27];
  assign T595 = T596 == T475;
  assign T596 = idxs[6'h28];
  assign T597 = {T600, T598};
  assign T598 = T599 == T475;
  assign T599 = idxs[6'h29];
  assign T600 = T601 == T475;
  assign T601 = idxs[6'h2a];
  assign T602 = {T608, T603};
  assign T603 = {T606, T604};
  assign T604 = T605 == T475;
  assign T605 = idxs[6'h2b];
  assign T606 = T607 == T475;
  assign T607 = idxs[6'h2c];
  assign T608 = {T611, T609};
  assign T609 = T610 == T475;
  assign T610 = idxs[6'h2d];
  assign T611 = T612 == T475;
  assign T612 = idxs[6'h2e];
  assign T613 = {T637, T614};
  assign T614 = {T626, T615};
  assign T615 = {T621, T616};
  assign T616 = {T619, T617};
  assign T617 = T618 == T475;
  assign T618 = idxs[6'h2f];
  assign T619 = T620 == T475;
  assign T620 = idxs[6'h30];
  assign T621 = {T624, T622};
  assign T622 = T623 == T475;
  assign T623 = idxs[6'h31];
  assign T624 = T625 == T475;
  assign T625 = idxs[6'h32];
  assign T626 = {T632, T627};
  assign T627 = {T630, T628};
  assign T628 = T629 == T475;
  assign T629 = idxs[6'h33];
  assign T630 = T631 == T475;
  assign T631 = idxs[6'h34];
  assign T632 = {T635, T633};
  assign T633 = T634 == T475;
  assign T634 = idxs[6'h35];
  assign T635 = T636 == T475;
  assign T636 = idxs[6'h36];
  assign T637 = {T649, T638};
  assign T638 = {T644, T639};
  assign T639 = {T642, T640};
  assign T640 = T641 == T475;
  assign T641 = idxs[6'h37];
  assign T642 = T643 == T475;
  assign T643 = idxs[6'h38];
  assign T644 = {T647, T645};
  assign T645 = T646 == T475;
  assign T646 = idxs[6'h39];
  assign T647 = T648 == T475;
  assign T648 = idxs[6'h3a];
  assign T649 = {T655, T650};
  assign T650 = {T653, T651};
  assign T651 = T652 == T475;
  assign T652 = idxs[6'h3b];
  assign T653 = T654 == T475;
  assign T654 = idxs[6'h3c];
  assign T655 = T656 == T475;
  assign T656 = idxs[6'h3d];
  assign T1607 = T1608[6'h3d:1'h0];
  assign T1608 = reset ? 64'h0 : T657;
  assign T657 = io_invalidate ? 64'h0 : T658;
  assign T658 = R7 ? T1038 : T1609;
  assign T1609 = {2'h0, T659};
  assign T659 = R7 ? T660 : idxValid;
  assign T660 = idxValid & T661;
  assign T661 = ~ T662;
  assign T662 = T663;
  assign T663 = {T853, T664};
  assign T664 = {T764, T665};
  assign T665 = {T717, T666};
  assign T666 = {T694, T667};
  assign T667 = {T683, T668};
  assign T668 = {T678, T669};
  assign T669 = T670 != 8'h0;
  assign T670 = pageReplEn & T1610;
  assign T1610 = {2'h0, T671};
  assign T671 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T672[3'h5:1'h0];
  assign T672 = 1'h1 << T673;
  assign T673 = tgtPages[6'h0];
  assign T1611 = {T1622, T1612};
  assign T1612 = {T1621, T1613};
  assign T1613 = T1614[1'h1:1'h1];
  assign T1614 = T1620 | T1615;
  assign T1615 = T1616[1'h1:1'h0];
  assign T1616 = T1619 | T1617;
  assign T1617 = T675[2'h3:1'h0];
  assign T675 = usePageHit ? T1618 : tgtPageRepl;
  assign T1618 = {2'h0, pageHit};
  assign T1619 = T675[3'h7:3'h4];
  assign T1620 = T1616[2'h3:2'h2];
  assign T1621 = T1620 != 2'h0;
  assign T1622 = T1619 != 4'h0;
  assign T676 = R7 & T677;
  assign T677 = T41 < 6'h3e;
  assign T678 = T679 != 8'h0;
  assign T679 = pageReplEn & T1623;
  assign T1623 = {2'h0, T680};
  assign T680 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T681[3'h5:1'h0];
  assign T681 = 1'h1 << T682;
  assign T682 = tgtPages[6'h1];
  assign T683 = {T689, T684};
  assign T684 = T685 != 8'h0;
  assign T685 = pageReplEn & T1624;
  assign T1624 = {2'h0, T686};
  assign T686 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T687[3'h5:1'h0];
  assign T687 = 1'h1 << T688;
  assign T688 = tgtPages[6'h2];
  assign T689 = T690 != 8'h0;
  assign T690 = pageReplEn & T1625;
  assign T1625 = {2'h0, T691};
  assign T691 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T692[3'h5:1'h0];
  assign T692 = 1'h1 << T693;
  assign T693 = tgtPages[6'h3];
  assign T694 = {T706, T695};
  assign T695 = {T701, T696};
  assign T696 = T697 != 8'h0;
  assign T697 = pageReplEn & T1626;
  assign T1626 = {2'h0, T698};
  assign T698 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T699[3'h5:1'h0];
  assign T699 = 1'h1 << T700;
  assign T700 = tgtPages[6'h4];
  assign T701 = T702 != 8'h0;
  assign T702 = pageReplEn & T1627;
  assign T1627 = {2'h0, T703};
  assign T703 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T704[3'h5:1'h0];
  assign T704 = 1'h1 << T705;
  assign T705 = tgtPages[6'h5];
  assign T706 = {T712, T707};
  assign T707 = T708 != 8'h0;
  assign T708 = pageReplEn & T1628;
  assign T1628 = {2'h0, T709};
  assign T709 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T710[3'h5:1'h0];
  assign T710 = 1'h1 << T711;
  assign T711 = tgtPages[6'h6];
  assign T712 = T713 != 8'h0;
  assign T713 = pageReplEn & T1629;
  assign T1629 = {2'h0, T714};
  assign T714 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T715[3'h5:1'h0];
  assign T715 = 1'h1 << T716;
  assign T716 = tgtPages[6'h7];
  assign T717 = {T741, T718};
  assign T718 = {T730, T719};
  assign T719 = {T725, T720};
  assign T720 = T721 != 8'h0;
  assign T721 = pageReplEn & T1630;
  assign T1630 = {2'h0, T722};
  assign T722 = idxPagesOH_8 | tgtPagesOH_8;
  assign tgtPagesOH_8 = T723[3'h5:1'h0];
  assign T723 = 1'h1 << T724;
  assign T724 = tgtPages[6'h8];
  assign T725 = T726 != 8'h0;
  assign T726 = pageReplEn & T1631;
  assign T1631 = {2'h0, T727};
  assign T727 = idxPagesOH_9 | tgtPagesOH_9;
  assign tgtPagesOH_9 = T728[3'h5:1'h0];
  assign T728 = 1'h1 << T729;
  assign T729 = tgtPages[6'h9];
  assign T730 = {T736, T731};
  assign T731 = T732 != 8'h0;
  assign T732 = pageReplEn & T1632;
  assign T1632 = {2'h0, T733};
  assign T733 = idxPagesOH_10 | tgtPagesOH_10;
  assign tgtPagesOH_10 = T734[3'h5:1'h0];
  assign T734 = 1'h1 << T735;
  assign T735 = tgtPages[6'ha];
  assign T736 = T737 != 8'h0;
  assign T737 = pageReplEn & T1633;
  assign T1633 = {2'h0, T738};
  assign T738 = idxPagesOH_11 | tgtPagesOH_11;
  assign tgtPagesOH_11 = T739[3'h5:1'h0];
  assign T739 = 1'h1 << T740;
  assign T740 = tgtPages[6'hb];
  assign T741 = {T753, T742};
  assign T742 = {T748, T743};
  assign T743 = T744 != 8'h0;
  assign T744 = pageReplEn & T1634;
  assign T1634 = {2'h0, T745};
  assign T745 = idxPagesOH_12 | tgtPagesOH_12;
  assign tgtPagesOH_12 = T746[3'h5:1'h0];
  assign T746 = 1'h1 << T747;
  assign T747 = tgtPages[6'hc];
  assign T748 = T749 != 8'h0;
  assign T749 = pageReplEn & T1635;
  assign T1635 = {2'h0, T750};
  assign T750 = idxPagesOH_13 | tgtPagesOH_13;
  assign tgtPagesOH_13 = T751[3'h5:1'h0];
  assign T751 = 1'h1 << T752;
  assign T752 = tgtPages[6'hd];
  assign T753 = {T759, T754};
  assign T754 = T755 != 8'h0;
  assign T755 = pageReplEn & T1636;
  assign T1636 = {2'h0, T756};
  assign T756 = idxPagesOH_14 | tgtPagesOH_14;
  assign tgtPagesOH_14 = T757[3'h5:1'h0];
  assign T757 = 1'h1 << T758;
  assign T758 = tgtPages[6'he];
  assign T759 = T760 != 8'h0;
  assign T760 = pageReplEn & T1637;
  assign T1637 = {2'h0, T761};
  assign T761 = idxPagesOH_15 | tgtPagesOH_15;
  assign tgtPagesOH_15 = T762[3'h5:1'h0];
  assign T762 = 1'h1 << T763;
  assign T763 = tgtPages[6'hf];
  assign T764 = {T812, T765};
  assign T765 = {T789, T766};
  assign T766 = {T778, T767};
  assign T767 = {T773, T768};
  assign T768 = T769 != 8'h0;
  assign T769 = pageReplEn & T1638;
  assign T1638 = {2'h0, T770};
  assign T770 = idxPagesOH_16 | tgtPagesOH_16;
  assign tgtPagesOH_16 = T771[3'h5:1'h0];
  assign T771 = 1'h1 << T772;
  assign T772 = tgtPages[6'h10];
  assign T773 = T774 != 8'h0;
  assign T774 = pageReplEn & T1639;
  assign T1639 = {2'h0, T775};
  assign T775 = idxPagesOH_17 | tgtPagesOH_17;
  assign tgtPagesOH_17 = T776[3'h5:1'h0];
  assign T776 = 1'h1 << T777;
  assign T777 = tgtPages[6'h11];
  assign T778 = {T784, T779};
  assign T779 = T780 != 8'h0;
  assign T780 = pageReplEn & T1640;
  assign T1640 = {2'h0, T781};
  assign T781 = idxPagesOH_18 | tgtPagesOH_18;
  assign tgtPagesOH_18 = T782[3'h5:1'h0];
  assign T782 = 1'h1 << T783;
  assign T783 = tgtPages[6'h12];
  assign T784 = T785 != 8'h0;
  assign T785 = pageReplEn & T1641;
  assign T1641 = {2'h0, T786};
  assign T786 = idxPagesOH_19 | tgtPagesOH_19;
  assign tgtPagesOH_19 = T787[3'h5:1'h0];
  assign T787 = 1'h1 << T788;
  assign T788 = tgtPages[6'h13];
  assign T789 = {T801, T790};
  assign T790 = {T796, T791};
  assign T791 = T792 != 8'h0;
  assign T792 = pageReplEn & T1642;
  assign T1642 = {2'h0, T793};
  assign T793 = idxPagesOH_20 | tgtPagesOH_20;
  assign tgtPagesOH_20 = T794[3'h5:1'h0];
  assign T794 = 1'h1 << T795;
  assign T795 = tgtPages[6'h14];
  assign T796 = T797 != 8'h0;
  assign T797 = pageReplEn & T1643;
  assign T1643 = {2'h0, T798};
  assign T798 = idxPagesOH_21 | tgtPagesOH_21;
  assign tgtPagesOH_21 = T799[3'h5:1'h0];
  assign T799 = 1'h1 << T800;
  assign T800 = tgtPages[6'h15];
  assign T801 = {T807, T802};
  assign T802 = T803 != 8'h0;
  assign T803 = pageReplEn & T1644;
  assign T1644 = {2'h0, T804};
  assign T804 = idxPagesOH_22 | tgtPagesOH_22;
  assign tgtPagesOH_22 = T805[3'h5:1'h0];
  assign T805 = 1'h1 << T806;
  assign T806 = tgtPages[6'h16];
  assign T807 = T808 != 8'h0;
  assign T808 = pageReplEn & T1645;
  assign T1645 = {2'h0, T809};
  assign T809 = idxPagesOH_23 | tgtPagesOH_23;
  assign tgtPagesOH_23 = T810[3'h5:1'h0];
  assign T810 = 1'h1 << T811;
  assign T811 = tgtPages[6'h17];
  assign T812 = {T836, T813};
  assign T813 = {T825, T814};
  assign T814 = {T820, T815};
  assign T815 = T816 != 8'h0;
  assign T816 = pageReplEn & T1646;
  assign T1646 = {2'h0, T817};
  assign T817 = idxPagesOH_24 | tgtPagesOH_24;
  assign tgtPagesOH_24 = T818[3'h5:1'h0];
  assign T818 = 1'h1 << T819;
  assign T819 = tgtPages[6'h18];
  assign T820 = T821 != 8'h0;
  assign T821 = pageReplEn & T1647;
  assign T1647 = {2'h0, T822};
  assign T822 = idxPagesOH_25 | tgtPagesOH_25;
  assign tgtPagesOH_25 = T823[3'h5:1'h0];
  assign T823 = 1'h1 << T824;
  assign T824 = tgtPages[6'h19];
  assign T825 = {T831, T826};
  assign T826 = T827 != 8'h0;
  assign T827 = pageReplEn & T1648;
  assign T1648 = {2'h0, T828};
  assign T828 = idxPagesOH_26 | tgtPagesOH_26;
  assign tgtPagesOH_26 = T829[3'h5:1'h0];
  assign T829 = 1'h1 << T830;
  assign T830 = tgtPages[6'h1a];
  assign T831 = T832 != 8'h0;
  assign T832 = pageReplEn & T1649;
  assign T1649 = {2'h0, T833};
  assign T833 = idxPagesOH_27 | tgtPagesOH_27;
  assign tgtPagesOH_27 = T834[3'h5:1'h0];
  assign T834 = 1'h1 << T835;
  assign T835 = tgtPages[6'h1b];
  assign T836 = {T848, T837};
  assign T837 = {T843, T838};
  assign T838 = T839 != 8'h0;
  assign T839 = pageReplEn & T1650;
  assign T1650 = {2'h0, T840};
  assign T840 = idxPagesOH_28 | tgtPagesOH_28;
  assign tgtPagesOH_28 = T841[3'h5:1'h0];
  assign T841 = 1'h1 << T842;
  assign T842 = tgtPages[6'h1c];
  assign T843 = T844 != 8'h0;
  assign T844 = pageReplEn & T1651;
  assign T1651 = {2'h0, T845};
  assign T845 = idxPagesOH_29 | tgtPagesOH_29;
  assign tgtPagesOH_29 = T846[3'h5:1'h0];
  assign T846 = 1'h1 << T847;
  assign T847 = tgtPages[6'h1d];
  assign T848 = T849 != 8'h0;
  assign T849 = pageReplEn & T1652;
  assign T1652 = {2'h0, T850};
  assign T850 = idxPagesOH_30 | tgtPagesOH_30;
  assign tgtPagesOH_30 = T851[3'h5:1'h0];
  assign T851 = 1'h1 << T852;
  assign T852 = tgtPages[6'h1e];
  assign T853 = {T949, T854};
  assign T854 = {T902, T855};
  assign T855 = {T879, T856};
  assign T856 = {T868, T857};
  assign T857 = {T863, T858};
  assign T858 = T859 != 8'h0;
  assign T859 = pageReplEn & T1653;
  assign T1653 = {2'h0, T860};
  assign T860 = idxPagesOH_31 | tgtPagesOH_31;
  assign tgtPagesOH_31 = T861[3'h5:1'h0];
  assign T861 = 1'h1 << T862;
  assign T862 = tgtPages[6'h1f];
  assign T863 = T864 != 8'h0;
  assign T864 = pageReplEn & T1654;
  assign T1654 = {2'h0, T865};
  assign T865 = idxPagesOH_32 | tgtPagesOH_32;
  assign tgtPagesOH_32 = T866[3'h5:1'h0];
  assign T866 = 1'h1 << T867;
  assign T867 = tgtPages[6'h20];
  assign T868 = {T874, T869};
  assign T869 = T870 != 8'h0;
  assign T870 = pageReplEn & T1655;
  assign T1655 = {2'h0, T871};
  assign T871 = idxPagesOH_33 | tgtPagesOH_33;
  assign tgtPagesOH_33 = T872[3'h5:1'h0];
  assign T872 = 1'h1 << T873;
  assign T873 = tgtPages[6'h21];
  assign T874 = T875 != 8'h0;
  assign T875 = pageReplEn & T1656;
  assign T1656 = {2'h0, T876};
  assign T876 = idxPagesOH_34 | tgtPagesOH_34;
  assign tgtPagesOH_34 = T877[3'h5:1'h0];
  assign T877 = 1'h1 << T878;
  assign T878 = tgtPages[6'h22];
  assign T879 = {T891, T880};
  assign T880 = {T886, T881};
  assign T881 = T882 != 8'h0;
  assign T882 = pageReplEn & T1657;
  assign T1657 = {2'h0, T883};
  assign T883 = idxPagesOH_35 | tgtPagesOH_35;
  assign tgtPagesOH_35 = T884[3'h5:1'h0];
  assign T884 = 1'h1 << T885;
  assign T885 = tgtPages[6'h23];
  assign T886 = T887 != 8'h0;
  assign T887 = pageReplEn & T1658;
  assign T1658 = {2'h0, T888};
  assign T888 = idxPagesOH_36 | tgtPagesOH_36;
  assign tgtPagesOH_36 = T889[3'h5:1'h0];
  assign T889 = 1'h1 << T890;
  assign T890 = tgtPages[6'h24];
  assign T891 = {T897, T892};
  assign T892 = T893 != 8'h0;
  assign T893 = pageReplEn & T1659;
  assign T1659 = {2'h0, T894};
  assign T894 = idxPagesOH_37 | tgtPagesOH_37;
  assign tgtPagesOH_37 = T895[3'h5:1'h0];
  assign T895 = 1'h1 << T896;
  assign T896 = tgtPages[6'h25];
  assign T897 = T898 != 8'h0;
  assign T898 = pageReplEn & T1660;
  assign T1660 = {2'h0, T899};
  assign T899 = idxPagesOH_38 | tgtPagesOH_38;
  assign tgtPagesOH_38 = T900[3'h5:1'h0];
  assign T900 = 1'h1 << T901;
  assign T901 = tgtPages[6'h26];
  assign T902 = {T926, T903};
  assign T903 = {T915, T904};
  assign T904 = {T910, T905};
  assign T905 = T906 != 8'h0;
  assign T906 = pageReplEn & T1661;
  assign T1661 = {2'h0, T907};
  assign T907 = idxPagesOH_39 | tgtPagesOH_39;
  assign tgtPagesOH_39 = T908[3'h5:1'h0];
  assign T908 = 1'h1 << T909;
  assign T909 = tgtPages[6'h27];
  assign T910 = T911 != 8'h0;
  assign T911 = pageReplEn & T1662;
  assign T1662 = {2'h0, T912};
  assign T912 = idxPagesOH_40 | tgtPagesOH_40;
  assign tgtPagesOH_40 = T913[3'h5:1'h0];
  assign T913 = 1'h1 << T914;
  assign T914 = tgtPages[6'h28];
  assign T915 = {T921, T916};
  assign T916 = T917 != 8'h0;
  assign T917 = pageReplEn & T1663;
  assign T1663 = {2'h0, T918};
  assign T918 = idxPagesOH_41 | tgtPagesOH_41;
  assign tgtPagesOH_41 = T919[3'h5:1'h0];
  assign T919 = 1'h1 << T920;
  assign T920 = tgtPages[6'h29];
  assign T921 = T922 != 8'h0;
  assign T922 = pageReplEn & T1664;
  assign T1664 = {2'h0, T923};
  assign T923 = idxPagesOH_42 | tgtPagesOH_42;
  assign tgtPagesOH_42 = T924[3'h5:1'h0];
  assign T924 = 1'h1 << T925;
  assign T925 = tgtPages[6'h2a];
  assign T926 = {T938, T927};
  assign T927 = {T933, T928};
  assign T928 = T929 != 8'h0;
  assign T929 = pageReplEn & T1665;
  assign T1665 = {2'h0, T930};
  assign T930 = idxPagesOH_43 | tgtPagesOH_43;
  assign tgtPagesOH_43 = T931[3'h5:1'h0];
  assign T931 = 1'h1 << T932;
  assign T932 = tgtPages[6'h2b];
  assign T933 = T934 != 8'h0;
  assign T934 = pageReplEn & T1666;
  assign T1666 = {2'h0, T935};
  assign T935 = idxPagesOH_44 | tgtPagesOH_44;
  assign tgtPagesOH_44 = T936[3'h5:1'h0];
  assign T936 = 1'h1 << T937;
  assign T937 = tgtPages[6'h2c];
  assign T938 = {T944, T939};
  assign T939 = T940 != 8'h0;
  assign T940 = pageReplEn & T1667;
  assign T1667 = {2'h0, T941};
  assign T941 = idxPagesOH_45 | tgtPagesOH_45;
  assign tgtPagesOH_45 = T942[3'h5:1'h0];
  assign T942 = 1'h1 << T943;
  assign T943 = tgtPages[6'h2d];
  assign T944 = T945 != 8'h0;
  assign T945 = pageReplEn & T1668;
  assign T1668 = {2'h0, T946};
  assign T946 = idxPagesOH_46 | tgtPagesOH_46;
  assign tgtPagesOH_46 = T947[3'h5:1'h0];
  assign T947 = 1'h1 << T948;
  assign T948 = tgtPages[6'h2e];
  assign T949 = {T997, T950};
  assign T950 = {T974, T951};
  assign T951 = {T963, T952};
  assign T952 = {T958, T953};
  assign T953 = T954 != 8'h0;
  assign T954 = pageReplEn & T1669;
  assign T1669 = {2'h0, T955};
  assign T955 = idxPagesOH_47 | tgtPagesOH_47;
  assign tgtPagesOH_47 = T956[3'h5:1'h0];
  assign T956 = 1'h1 << T957;
  assign T957 = tgtPages[6'h2f];
  assign T958 = T959 != 8'h0;
  assign T959 = pageReplEn & T1670;
  assign T1670 = {2'h0, T960};
  assign T960 = idxPagesOH_48 | tgtPagesOH_48;
  assign tgtPagesOH_48 = T961[3'h5:1'h0];
  assign T961 = 1'h1 << T962;
  assign T962 = tgtPages[6'h30];
  assign T963 = {T969, T964};
  assign T964 = T965 != 8'h0;
  assign T965 = pageReplEn & T1671;
  assign T1671 = {2'h0, T966};
  assign T966 = idxPagesOH_49 | tgtPagesOH_49;
  assign tgtPagesOH_49 = T967[3'h5:1'h0];
  assign T967 = 1'h1 << T968;
  assign T968 = tgtPages[6'h31];
  assign T969 = T970 != 8'h0;
  assign T970 = pageReplEn & T1672;
  assign T1672 = {2'h0, T971};
  assign T971 = idxPagesOH_50 | tgtPagesOH_50;
  assign tgtPagesOH_50 = T972[3'h5:1'h0];
  assign T972 = 1'h1 << T973;
  assign T973 = tgtPages[6'h32];
  assign T974 = {T986, T975};
  assign T975 = {T981, T976};
  assign T976 = T977 != 8'h0;
  assign T977 = pageReplEn & T1673;
  assign T1673 = {2'h0, T978};
  assign T978 = idxPagesOH_51 | tgtPagesOH_51;
  assign tgtPagesOH_51 = T979[3'h5:1'h0];
  assign T979 = 1'h1 << T980;
  assign T980 = tgtPages[6'h33];
  assign T981 = T982 != 8'h0;
  assign T982 = pageReplEn & T1674;
  assign T1674 = {2'h0, T983};
  assign T983 = idxPagesOH_52 | tgtPagesOH_52;
  assign tgtPagesOH_52 = T984[3'h5:1'h0];
  assign T984 = 1'h1 << T985;
  assign T985 = tgtPages[6'h34];
  assign T986 = {T992, T987};
  assign T987 = T988 != 8'h0;
  assign T988 = pageReplEn & T1675;
  assign T1675 = {2'h0, T989};
  assign T989 = idxPagesOH_53 | tgtPagesOH_53;
  assign tgtPagesOH_53 = T990[3'h5:1'h0];
  assign T990 = 1'h1 << T991;
  assign T991 = tgtPages[6'h35];
  assign T992 = T993 != 8'h0;
  assign T993 = pageReplEn & T1676;
  assign T1676 = {2'h0, T994};
  assign T994 = idxPagesOH_54 | tgtPagesOH_54;
  assign tgtPagesOH_54 = T995[3'h5:1'h0];
  assign T995 = 1'h1 << T996;
  assign T996 = tgtPages[6'h36];
  assign T997 = {T1021, T998};
  assign T998 = {T1010, T999};
  assign T999 = {T1005, T1000};
  assign T1000 = T1001 != 8'h0;
  assign T1001 = pageReplEn & T1677;
  assign T1677 = {2'h0, T1002};
  assign T1002 = idxPagesOH_55 | tgtPagesOH_55;
  assign tgtPagesOH_55 = T1003[3'h5:1'h0];
  assign T1003 = 1'h1 << T1004;
  assign T1004 = tgtPages[6'h37];
  assign T1005 = T1006 != 8'h0;
  assign T1006 = pageReplEn & T1678;
  assign T1678 = {2'h0, T1007};
  assign T1007 = idxPagesOH_56 | tgtPagesOH_56;
  assign tgtPagesOH_56 = T1008[3'h5:1'h0];
  assign T1008 = 1'h1 << T1009;
  assign T1009 = tgtPages[6'h38];
  assign T1010 = {T1016, T1011};
  assign T1011 = T1012 != 8'h0;
  assign T1012 = pageReplEn & T1679;
  assign T1679 = {2'h0, T1013};
  assign T1013 = idxPagesOH_57 | tgtPagesOH_57;
  assign tgtPagesOH_57 = T1014[3'h5:1'h0];
  assign T1014 = 1'h1 << T1015;
  assign T1015 = tgtPages[6'h39];
  assign T1016 = T1017 != 8'h0;
  assign T1017 = pageReplEn & T1680;
  assign T1680 = {2'h0, T1018};
  assign T1018 = idxPagesOH_58 | tgtPagesOH_58;
  assign tgtPagesOH_58 = T1019[3'h5:1'h0];
  assign T1019 = 1'h1 << T1020;
  assign T1020 = tgtPages[6'h3a];
  assign T1021 = {T1033, T1022};
  assign T1022 = {T1028, T1023};
  assign T1023 = T1024 != 8'h0;
  assign T1024 = pageReplEn & T1681;
  assign T1681 = {2'h0, T1025};
  assign T1025 = idxPagesOH_59 | tgtPagesOH_59;
  assign tgtPagesOH_59 = T1026[3'h5:1'h0];
  assign T1026 = 1'h1 << T1027;
  assign T1027 = tgtPages[6'h3b];
  assign T1028 = T1029 != 8'h0;
  assign T1029 = pageReplEn & T1682;
  assign T1682 = {2'h0, T1030};
  assign T1030 = idxPagesOH_60 | tgtPagesOH_60;
  assign tgtPagesOH_60 = T1031[3'h5:1'h0];
  assign T1031 = 1'h1 << T1032;
  assign T1032 = tgtPages[6'h3c];
  assign T1033 = T1034 != 8'h0;
  assign T1034 = pageReplEn & T1683;
  assign T1683 = {2'h0, T1035};
  assign T1035 = idxPagesOH_61 | tgtPagesOH_61;
  assign tgtPagesOH_61 = T1036[3'h5:1'h0];
  assign T1036 = 1'h1 << T1037;
  assign T1037 = tgtPages[6'h3d];
  assign T1038 = T1045 | T1039;
  assign T1039 = T1685 & T1040;
  assign T1040 = T1042 | T1684;
  assign T1684 = {2'h0, T1041};
  assign T1041 = idxValid ^ idxValid;
  assign T1042 = 1'h1 << T41;
  assign T1685 = T1043 ? 64'hffffffffffffffff : 64'h0;
  assign T1043 = T1044;
  assign T1044 = 1'h1;
  assign T1045 = T1686 & T1046;
  assign T1046 = ~ T1040;
  assign T1686 = {2'h0, T659};
  assign T1047 = io_req_valid & T1048;
  assign T1048 = hits != 62'h0;
  assign T1049 = {io_bht_update_bits_taken, T1050};
  assign T1050 = io_bht_update_bits_prediction_bits_bht_history[3'h6:1'h1];
  assign T1051 = T21 & io_bht_update_bits_mispredict;
  assign T1052 = io_req_bits_addr[4'h8:2'h2];
  assign io_resp_bits_bht_history = T1053;
  assign T1053 = R25;
  assign io_resp_bits_entry = T1687;
  assign T1687 = {T1712, T1688};
  assign T1688 = {T1711, T1689};
  assign T1689 = {T1710, T1690};
  assign T1690 = {T1709, T1691};
  assign T1691 = {T1708, T1692};
  assign T1692 = T1693[1'h1:1'h1];
  assign T1693 = T1707 | T1694;
  assign T1694 = T1695[1'h1:1'h0];
  assign T1695 = T1706 | T1696;
  assign T1696 = T1697[2'h3:1'h0];
  assign T1697 = T1705 | T1698;
  assign T1698 = T1699[3'h7:1'h0];
  assign T1699 = T1704 | T1700;
  assign T1700 = T1701[4'hf:1'h0];
  assign T1701 = T1703 | T1702;
  assign T1702 = hits[5'h1f:1'h0];
  assign T1703 = hits[6'h3d:6'h20];
  assign T1704 = T1701[5'h1f:5'h10];
  assign T1705 = T1699[4'hf:4'h8];
  assign T1706 = T1697[3'h7:3'h4];
  assign T1707 = T1695[2'h3:2'h2];
  assign T1708 = T1707 != 2'h0;
  assign T1709 = T1706 != 4'h0;
  assign T1710 = T1705 != 8'h0;
  assign T1711 = T1704 != 16'h0;
  assign T1712 = T1703 != 30'h0;
  assign io_resp_bits_target = T1055;
  assign T1055 = T1566 ? io_ras_update_bits_returnAddr : T1056;
  assign T1056 = T1549 ? T1516 : T1057;
  assign T1057 = {T1308, T1058};
  assign T1058 = T1065 | T1059;
  assign T1059 = T1064 ? T1060 : 13'h0;
  assign T1060 = tgts[6'h3d];
  assign T1713 = io_req_bits_addr[4'hc:1'h0];
  assign T1062 = R7 & T1063;
  assign T1063 = T41 < 6'h3e;
  assign T1064 = hits[6'h3d:6'h3d];
  assign T1065 = T1069 | T1066;
  assign T1066 = T1068 ? T1067 : 13'h0;
  assign T1067 = tgts[6'h3c];
  assign T1068 = hits[6'h3c:6'h3c];
  assign T1069 = T1073 | T1070;
  assign T1070 = T1072 ? T1071 : 13'h0;
  assign T1071 = tgts[6'h3b];
  assign T1072 = hits[6'h3b:6'h3b];
  assign T1073 = T1077 | T1074;
  assign T1074 = T1076 ? T1075 : 13'h0;
  assign T1075 = tgts[6'h3a];
  assign T1076 = hits[6'h3a:6'h3a];
  assign T1077 = T1081 | T1078;
  assign T1078 = T1080 ? T1079 : 13'h0;
  assign T1079 = tgts[6'h39];
  assign T1080 = hits[6'h39:6'h39];
  assign T1081 = T1085 | T1082;
  assign T1082 = T1084 ? T1083 : 13'h0;
  assign T1083 = tgts[6'h38];
  assign T1084 = hits[6'h38:6'h38];
  assign T1085 = T1089 | T1086;
  assign T1086 = T1088 ? T1087 : 13'h0;
  assign T1087 = tgts[6'h37];
  assign T1088 = hits[6'h37:6'h37];
  assign T1089 = T1093 | T1090;
  assign T1090 = T1092 ? T1091 : 13'h0;
  assign T1091 = tgts[6'h36];
  assign T1092 = hits[6'h36:6'h36];
  assign T1093 = T1097 | T1094;
  assign T1094 = T1096 ? T1095 : 13'h0;
  assign T1095 = tgts[6'h35];
  assign T1096 = hits[6'h35:6'h35];
  assign T1097 = T1101 | T1098;
  assign T1098 = T1100 ? T1099 : 13'h0;
  assign T1099 = tgts[6'h34];
  assign T1100 = hits[6'h34:6'h34];
  assign T1101 = T1105 | T1102;
  assign T1102 = T1104 ? T1103 : 13'h0;
  assign T1103 = tgts[6'h33];
  assign T1104 = hits[6'h33:6'h33];
  assign T1105 = T1109 | T1106;
  assign T1106 = T1108 ? T1107 : 13'h0;
  assign T1107 = tgts[6'h32];
  assign T1108 = hits[6'h32:6'h32];
  assign T1109 = T1113 | T1110;
  assign T1110 = T1112 ? T1111 : 13'h0;
  assign T1111 = tgts[6'h31];
  assign T1112 = hits[6'h31:6'h31];
  assign T1113 = T1117 | T1114;
  assign T1114 = T1116 ? T1115 : 13'h0;
  assign T1115 = tgts[6'h30];
  assign T1116 = hits[6'h30:6'h30];
  assign T1117 = T1121 | T1118;
  assign T1118 = T1120 ? T1119 : 13'h0;
  assign T1119 = tgts[6'h2f];
  assign T1120 = hits[6'h2f:6'h2f];
  assign T1121 = T1125 | T1122;
  assign T1122 = T1124 ? T1123 : 13'h0;
  assign T1123 = tgts[6'h2e];
  assign T1124 = hits[6'h2e:6'h2e];
  assign T1125 = T1129 | T1126;
  assign T1126 = T1128 ? T1127 : 13'h0;
  assign T1127 = tgts[6'h2d];
  assign T1128 = hits[6'h2d:6'h2d];
  assign T1129 = T1133 | T1130;
  assign T1130 = T1132 ? T1131 : 13'h0;
  assign T1131 = tgts[6'h2c];
  assign T1132 = hits[6'h2c:6'h2c];
  assign T1133 = T1137 | T1134;
  assign T1134 = T1136 ? T1135 : 13'h0;
  assign T1135 = tgts[6'h2b];
  assign T1136 = hits[6'h2b:6'h2b];
  assign T1137 = T1141 | T1138;
  assign T1138 = T1140 ? T1139 : 13'h0;
  assign T1139 = tgts[6'h2a];
  assign T1140 = hits[6'h2a:6'h2a];
  assign T1141 = T1145 | T1142;
  assign T1142 = T1144 ? T1143 : 13'h0;
  assign T1143 = tgts[6'h29];
  assign T1144 = hits[6'h29:6'h29];
  assign T1145 = T1149 | T1146;
  assign T1146 = T1148 ? T1147 : 13'h0;
  assign T1147 = tgts[6'h28];
  assign T1148 = hits[6'h28:6'h28];
  assign T1149 = T1153 | T1150;
  assign T1150 = T1152 ? T1151 : 13'h0;
  assign T1151 = tgts[6'h27];
  assign T1152 = hits[6'h27:6'h27];
  assign T1153 = T1157 | T1154;
  assign T1154 = T1156 ? T1155 : 13'h0;
  assign T1155 = tgts[6'h26];
  assign T1156 = hits[6'h26:6'h26];
  assign T1157 = T1161 | T1158;
  assign T1158 = T1160 ? T1159 : 13'h0;
  assign T1159 = tgts[6'h25];
  assign T1160 = hits[6'h25:6'h25];
  assign T1161 = T1165 | T1162;
  assign T1162 = T1164 ? T1163 : 13'h0;
  assign T1163 = tgts[6'h24];
  assign T1164 = hits[6'h24:6'h24];
  assign T1165 = T1169 | T1166;
  assign T1166 = T1168 ? T1167 : 13'h0;
  assign T1167 = tgts[6'h23];
  assign T1168 = hits[6'h23:6'h23];
  assign T1169 = T1173 | T1170;
  assign T1170 = T1172 ? T1171 : 13'h0;
  assign T1171 = tgts[6'h22];
  assign T1172 = hits[6'h22:6'h22];
  assign T1173 = T1177 | T1174;
  assign T1174 = T1176 ? T1175 : 13'h0;
  assign T1175 = tgts[6'h21];
  assign T1176 = hits[6'h21:6'h21];
  assign T1177 = T1181 | T1178;
  assign T1178 = T1180 ? T1179 : 13'h0;
  assign T1179 = tgts[6'h20];
  assign T1180 = hits[6'h20:6'h20];
  assign T1181 = T1185 | T1182;
  assign T1182 = T1184 ? T1183 : 13'h0;
  assign T1183 = tgts[6'h1f];
  assign T1184 = hits[5'h1f:5'h1f];
  assign T1185 = T1189 | T1186;
  assign T1186 = T1188 ? T1187 : 13'h0;
  assign T1187 = tgts[6'h1e];
  assign T1188 = hits[5'h1e:5'h1e];
  assign T1189 = T1193 | T1190;
  assign T1190 = T1192 ? T1191 : 13'h0;
  assign T1191 = tgts[6'h1d];
  assign T1192 = hits[5'h1d:5'h1d];
  assign T1193 = T1197 | T1194;
  assign T1194 = T1196 ? T1195 : 13'h0;
  assign T1195 = tgts[6'h1c];
  assign T1196 = hits[5'h1c:5'h1c];
  assign T1197 = T1201 | T1198;
  assign T1198 = T1200 ? T1199 : 13'h0;
  assign T1199 = tgts[6'h1b];
  assign T1200 = hits[5'h1b:5'h1b];
  assign T1201 = T1205 | T1202;
  assign T1202 = T1204 ? T1203 : 13'h0;
  assign T1203 = tgts[6'h1a];
  assign T1204 = hits[5'h1a:5'h1a];
  assign T1205 = T1209 | T1206;
  assign T1206 = T1208 ? T1207 : 13'h0;
  assign T1207 = tgts[6'h19];
  assign T1208 = hits[5'h19:5'h19];
  assign T1209 = T1213 | T1210;
  assign T1210 = T1212 ? T1211 : 13'h0;
  assign T1211 = tgts[6'h18];
  assign T1212 = hits[5'h18:5'h18];
  assign T1213 = T1217 | T1214;
  assign T1214 = T1216 ? T1215 : 13'h0;
  assign T1215 = tgts[6'h17];
  assign T1216 = hits[5'h17:5'h17];
  assign T1217 = T1221 | T1218;
  assign T1218 = T1220 ? T1219 : 13'h0;
  assign T1219 = tgts[6'h16];
  assign T1220 = hits[5'h16:5'h16];
  assign T1221 = T1225 | T1222;
  assign T1222 = T1224 ? T1223 : 13'h0;
  assign T1223 = tgts[6'h15];
  assign T1224 = hits[5'h15:5'h15];
  assign T1225 = T1229 | T1226;
  assign T1226 = T1228 ? T1227 : 13'h0;
  assign T1227 = tgts[6'h14];
  assign T1228 = hits[5'h14:5'h14];
  assign T1229 = T1233 | T1230;
  assign T1230 = T1232 ? T1231 : 13'h0;
  assign T1231 = tgts[6'h13];
  assign T1232 = hits[5'h13:5'h13];
  assign T1233 = T1237 | T1234;
  assign T1234 = T1236 ? T1235 : 13'h0;
  assign T1235 = tgts[6'h12];
  assign T1236 = hits[5'h12:5'h12];
  assign T1237 = T1241 | T1238;
  assign T1238 = T1240 ? T1239 : 13'h0;
  assign T1239 = tgts[6'h11];
  assign T1240 = hits[5'h11:5'h11];
  assign T1241 = T1245 | T1242;
  assign T1242 = T1244 ? T1243 : 13'h0;
  assign T1243 = tgts[6'h10];
  assign T1244 = hits[5'h10:5'h10];
  assign T1245 = T1249 | T1246;
  assign T1246 = T1248 ? T1247 : 13'h0;
  assign T1247 = tgts[6'hf];
  assign T1248 = hits[4'hf:4'hf];
  assign T1249 = T1253 | T1250;
  assign T1250 = T1252 ? T1251 : 13'h0;
  assign T1251 = tgts[6'he];
  assign T1252 = hits[4'he:4'he];
  assign T1253 = T1257 | T1254;
  assign T1254 = T1256 ? T1255 : 13'h0;
  assign T1255 = tgts[6'hd];
  assign T1256 = hits[4'hd:4'hd];
  assign T1257 = T1261 | T1258;
  assign T1258 = T1260 ? T1259 : 13'h0;
  assign T1259 = tgts[6'hc];
  assign T1260 = hits[4'hc:4'hc];
  assign T1261 = T1265 | T1262;
  assign T1262 = T1264 ? T1263 : 13'h0;
  assign T1263 = tgts[6'hb];
  assign T1264 = hits[4'hb:4'hb];
  assign T1265 = T1269 | T1266;
  assign T1266 = T1268 ? T1267 : 13'h0;
  assign T1267 = tgts[6'ha];
  assign T1268 = hits[4'ha:4'ha];
  assign T1269 = T1273 | T1270;
  assign T1270 = T1272 ? T1271 : 13'h0;
  assign T1271 = tgts[6'h9];
  assign T1272 = hits[4'h9:4'h9];
  assign T1273 = T1277 | T1274;
  assign T1274 = T1276 ? T1275 : 13'h0;
  assign T1275 = tgts[6'h8];
  assign T1276 = hits[4'h8:4'h8];
  assign T1277 = T1281 | T1278;
  assign T1278 = T1280 ? T1279 : 13'h0;
  assign T1279 = tgts[6'h7];
  assign T1280 = hits[3'h7:3'h7];
  assign T1281 = T1285 | T1282;
  assign T1282 = T1284 ? T1283 : 13'h0;
  assign T1283 = tgts[6'h6];
  assign T1284 = hits[3'h6:3'h6];
  assign T1285 = T1289 | T1286;
  assign T1286 = T1288 ? T1287 : 13'h0;
  assign T1287 = tgts[6'h5];
  assign T1288 = hits[3'h5:3'h5];
  assign T1289 = T1293 | T1290;
  assign T1290 = T1292 ? T1291 : 13'h0;
  assign T1291 = tgts[6'h4];
  assign T1292 = hits[3'h4:3'h4];
  assign T1293 = T1297 | T1294;
  assign T1294 = T1296 ? T1295 : 13'h0;
  assign T1295 = tgts[6'h3];
  assign T1296 = hits[2'h3:2'h3];
  assign T1297 = T1301 | T1298;
  assign T1298 = T1300 ? T1299 : 13'h0;
  assign T1299 = tgts[6'h2];
  assign T1300 = hits[2'h2:2'h2];
  assign T1301 = T1305 | T1302;
  assign T1302 = T1304 ? T1303 : 13'h0;
  assign T1303 = tgts[6'h1];
  assign T1304 = hits[1'h1:1'h1];
  assign T1305 = T1307 ? T1306 : 13'h0;
  assign T1306 = tgts[6'h0];
  assign T1307 = hits[1'h0:1'h0];
  assign T1308 = T1497 | T1309;
  assign T1309 = T1311 ? T1310 : 30'h0;
  assign T1310 = pages[3'h5];
  assign T1311 = T1312[3'h5:3'h5];
  assign T1312 = T1315 | T1313;
  assign T1313 = T1314 ? tgtPagesOH_61 : 6'h0;
  assign T1314 = hits[6'h3d:6'h3d];
  assign T1315 = T1318 | T1316;
  assign T1316 = T1317 ? tgtPagesOH_60 : 6'h0;
  assign T1317 = hits[6'h3c:6'h3c];
  assign T1318 = T1321 | T1319;
  assign T1319 = T1320 ? tgtPagesOH_59 : 6'h0;
  assign T1320 = hits[6'h3b:6'h3b];
  assign T1321 = T1324 | T1322;
  assign T1322 = T1323 ? tgtPagesOH_58 : 6'h0;
  assign T1323 = hits[6'h3a:6'h3a];
  assign T1324 = T1327 | T1325;
  assign T1325 = T1326 ? tgtPagesOH_57 : 6'h0;
  assign T1326 = hits[6'h39:6'h39];
  assign T1327 = T1330 | T1328;
  assign T1328 = T1329 ? tgtPagesOH_56 : 6'h0;
  assign T1329 = hits[6'h38:6'h38];
  assign T1330 = T1333 | T1331;
  assign T1331 = T1332 ? tgtPagesOH_55 : 6'h0;
  assign T1332 = hits[6'h37:6'h37];
  assign T1333 = T1336 | T1334;
  assign T1334 = T1335 ? tgtPagesOH_54 : 6'h0;
  assign T1335 = hits[6'h36:6'h36];
  assign T1336 = T1339 | T1337;
  assign T1337 = T1338 ? tgtPagesOH_53 : 6'h0;
  assign T1338 = hits[6'h35:6'h35];
  assign T1339 = T1342 | T1340;
  assign T1340 = T1341 ? tgtPagesOH_52 : 6'h0;
  assign T1341 = hits[6'h34:6'h34];
  assign T1342 = T1345 | T1343;
  assign T1343 = T1344 ? tgtPagesOH_51 : 6'h0;
  assign T1344 = hits[6'h33:6'h33];
  assign T1345 = T1348 | T1346;
  assign T1346 = T1347 ? tgtPagesOH_50 : 6'h0;
  assign T1347 = hits[6'h32:6'h32];
  assign T1348 = T1351 | T1349;
  assign T1349 = T1350 ? tgtPagesOH_49 : 6'h0;
  assign T1350 = hits[6'h31:6'h31];
  assign T1351 = T1354 | T1352;
  assign T1352 = T1353 ? tgtPagesOH_48 : 6'h0;
  assign T1353 = hits[6'h30:6'h30];
  assign T1354 = T1357 | T1355;
  assign T1355 = T1356 ? tgtPagesOH_47 : 6'h0;
  assign T1356 = hits[6'h2f:6'h2f];
  assign T1357 = T1360 | T1358;
  assign T1358 = T1359 ? tgtPagesOH_46 : 6'h0;
  assign T1359 = hits[6'h2e:6'h2e];
  assign T1360 = T1363 | T1361;
  assign T1361 = T1362 ? tgtPagesOH_45 : 6'h0;
  assign T1362 = hits[6'h2d:6'h2d];
  assign T1363 = T1366 | T1364;
  assign T1364 = T1365 ? tgtPagesOH_44 : 6'h0;
  assign T1365 = hits[6'h2c:6'h2c];
  assign T1366 = T1369 | T1367;
  assign T1367 = T1368 ? tgtPagesOH_43 : 6'h0;
  assign T1368 = hits[6'h2b:6'h2b];
  assign T1369 = T1372 | T1370;
  assign T1370 = T1371 ? tgtPagesOH_42 : 6'h0;
  assign T1371 = hits[6'h2a:6'h2a];
  assign T1372 = T1375 | T1373;
  assign T1373 = T1374 ? tgtPagesOH_41 : 6'h0;
  assign T1374 = hits[6'h29:6'h29];
  assign T1375 = T1378 | T1376;
  assign T1376 = T1377 ? tgtPagesOH_40 : 6'h0;
  assign T1377 = hits[6'h28:6'h28];
  assign T1378 = T1381 | T1379;
  assign T1379 = T1380 ? tgtPagesOH_39 : 6'h0;
  assign T1380 = hits[6'h27:6'h27];
  assign T1381 = T1384 | T1382;
  assign T1382 = T1383 ? tgtPagesOH_38 : 6'h0;
  assign T1383 = hits[6'h26:6'h26];
  assign T1384 = T1387 | T1385;
  assign T1385 = T1386 ? tgtPagesOH_37 : 6'h0;
  assign T1386 = hits[6'h25:6'h25];
  assign T1387 = T1390 | T1388;
  assign T1388 = T1389 ? tgtPagesOH_36 : 6'h0;
  assign T1389 = hits[6'h24:6'h24];
  assign T1390 = T1393 | T1391;
  assign T1391 = T1392 ? tgtPagesOH_35 : 6'h0;
  assign T1392 = hits[6'h23:6'h23];
  assign T1393 = T1396 | T1394;
  assign T1394 = T1395 ? tgtPagesOH_34 : 6'h0;
  assign T1395 = hits[6'h22:6'h22];
  assign T1396 = T1399 | T1397;
  assign T1397 = T1398 ? tgtPagesOH_33 : 6'h0;
  assign T1398 = hits[6'h21:6'h21];
  assign T1399 = T1402 | T1400;
  assign T1400 = T1401 ? tgtPagesOH_32 : 6'h0;
  assign T1401 = hits[6'h20:6'h20];
  assign T1402 = T1405 | T1403;
  assign T1403 = T1404 ? tgtPagesOH_31 : 6'h0;
  assign T1404 = hits[5'h1f:5'h1f];
  assign T1405 = T1408 | T1406;
  assign T1406 = T1407 ? tgtPagesOH_30 : 6'h0;
  assign T1407 = hits[5'h1e:5'h1e];
  assign T1408 = T1411 | T1409;
  assign T1409 = T1410 ? tgtPagesOH_29 : 6'h0;
  assign T1410 = hits[5'h1d:5'h1d];
  assign T1411 = T1414 | T1412;
  assign T1412 = T1413 ? tgtPagesOH_28 : 6'h0;
  assign T1413 = hits[5'h1c:5'h1c];
  assign T1414 = T1417 | T1415;
  assign T1415 = T1416 ? tgtPagesOH_27 : 6'h0;
  assign T1416 = hits[5'h1b:5'h1b];
  assign T1417 = T1420 | T1418;
  assign T1418 = T1419 ? tgtPagesOH_26 : 6'h0;
  assign T1419 = hits[5'h1a:5'h1a];
  assign T1420 = T1423 | T1421;
  assign T1421 = T1422 ? tgtPagesOH_25 : 6'h0;
  assign T1422 = hits[5'h19:5'h19];
  assign T1423 = T1426 | T1424;
  assign T1424 = T1425 ? tgtPagesOH_24 : 6'h0;
  assign T1425 = hits[5'h18:5'h18];
  assign T1426 = T1429 | T1427;
  assign T1427 = T1428 ? tgtPagesOH_23 : 6'h0;
  assign T1428 = hits[5'h17:5'h17];
  assign T1429 = T1432 | T1430;
  assign T1430 = T1431 ? tgtPagesOH_22 : 6'h0;
  assign T1431 = hits[5'h16:5'h16];
  assign T1432 = T1435 | T1433;
  assign T1433 = T1434 ? tgtPagesOH_21 : 6'h0;
  assign T1434 = hits[5'h15:5'h15];
  assign T1435 = T1438 | T1436;
  assign T1436 = T1437 ? tgtPagesOH_20 : 6'h0;
  assign T1437 = hits[5'h14:5'h14];
  assign T1438 = T1441 | T1439;
  assign T1439 = T1440 ? tgtPagesOH_19 : 6'h0;
  assign T1440 = hits[5'h13:5'h13];
  assign T1441 = T1444 | T1442;
  assign T1442 = T1443 ? tgtPagesOH_18 : 6'h0;
  assign T1443 = hits[5'h12:5'h12];
  assign T1444 = T1447 | T1445;
  assign T1445 = T1446 ? tgtPagesOH_17 : 6'h0;
  assign T1446 = hits[5'h11:5'h11];
  assign T1447 = T1450 | T1448;
  assign T1448 = T1449 ? tgtPagesOH_16 : 6'h0;
  assign T1449 = hits[5'h10:5'h10];
  assign T1450 = T1453 | T1451;
  assign T1451 = T1452 ? tgtPagesOH_15 : 6'h0;
  assign T1452 = hits[4'hf:4'hf];
  assign T1453 = T1456 | T1454;
  assign T1454 = T1455 ? tgtPagesOH_14 : 6'h0;
  assign T1455 = hits[4'he:4'he];
  assign T1456 = T1459 | T1457;
  assign T1457 = T1458 ? tgtPagesOH_13 : 6'h0;
  assign T1458 = hits[4'hd:4'hd];
  assign T1459 = T1462 | T1460;
  assign T1460 = T1461 ? tgtPagesOH_12 : 6'h0;
  assign T1461 = hits[4'hc:4'hc];
  assign T1462 = T1465 | T1463;
  assign T1463 = T1464 ? tgtPagesOH_11 : 6'h0;
  assign T1464 = hits[4'hb:4'hb];
  assign T1465 = T1468 | T1466;
  assign T1466 = T1467 ? tgtPagesOH_10 : 6'h0;
  assign T1467 = hits[4'ha:4'ha];
  assign T1468 = T1471 | T1469;
  assign T1469 = T1470 ? tgtPagesOH_9 : 6'h0;
  assign T1470 = hits[4'h9:4'h9];
  assign T1471 = T1474 | T1472;
  assign T1472 = T1473 ? tgtPagesOH_8 : 6'h0;
  assign T1473 = hits[4'h8:4'h8];
  assign T1474 = T1477 | T1475;
  assign T1475 = T1476 ? tgtPagesOH_7 : 6'h0;
  assign T1476 = hits[3'h7:3'h7];
  assign T1477 = T1480 | T1478;
  assign T1478 = T1479 ? tgtPagesOH_6 : 6'h0;
  assign T1479 = hits[3'h6:3'h6];
  assign T1480 = T1483 | T1481;
  assign T1481 = T1482 ? tgtPagesOH_5 : 6'h0;
  assign T1482 = hits[3'h5:3'h5];
  assign T1483 = T1486 | T1484;
  assign T1484 = T1485 ? tgtPagesOH_4 : 6'h0;
  assign T1485 = hits[3'h4:3'h4];
  assign T1486 = T1489 | T1487;
  assign T1487 = T1488 ? tgtPagesOH_3 : 6'h0;
  assign T1488 = hits[2'h3:2'h3];
  assign T1489 = T1492 | T1490;
  assign T1490 = T1491 ? tgtPagesOH_2 : 6'h0;
  assign T1491 = hits[2'h2:2'h2];
  assign T1492 = T1495 | T1493;
  assign T1493 = T1494 ? tgtPagesOH_1 : 6'h0;
  assign T1494 = hits[1'h1:1'h1];
  assign T1495 = T1496 ? tgtPagesOH_0 : 6'h0;
  assign T1496 = hits[1'h0:1'h0];
  assign T1497 = T1501 | T1498;
  assign T1498 = T1500 ? T1499 : 30'h0;
  assign T1499 = pages[3'h4];
  assign T1500 = T1312[3'h4:3'h4];
  assign T1501 = T1505 | T1502;
  assign T1502 = T1504 ? T1503 : 30'h0;
  assign T1503 = pages[3'h3];
  assign T1504 = T1312[2'h3:2'h3];
  assign T1505 = T1509 | T1506;
  assign T1506 = T1508 ? T1507 : 30'h0;
  assign T1507 = pages[3'h2];
  assign T1508 = T1312[2'h2:2'h2];
  assign T1509 = T1513 | T1510;
  assign T1510 = T1512 ? T1511 : 30'h0;
  assign T1511 = pages[3'h1];
  assign T1512 = T1312[1'h1:1'h1];
  assign T1513 = T1515 ? T1514 : 30'h0;
  assign T1514 = pages[3'h0];
  assign T1515 = T1312[1'h0:1'h0];
  assign T1516 = T1548 ? R1544 : R1517;
  assign T1518 = T1519 ? io_ras_update_bits_returnAddr : R1517;
  assign T1519 = T1543 & T1520;
  assign T1520 = T1521[1'h0:1'h0];
  assign T1521 = 1'h1 << T1522;
  assign T1522 = T1523;
  assign T1523 = R1524 + 1'h1;
  assign T1714 = reset ? 1'h0 : T1525;
  assign T1525 = T1528 ? T1527 : T1526;
  assign T1526 = T1543 ? T1523 : R1524;
  assign T1527 = R1524 - 1'h1;
  assign T1528 = T1539 & T1529;
  assign T1529 = T1530 ^ 1'h1;
  assign T1530 = R1531 == 2'h0;
  assign T1715 = reset ? 2'h0 : T1532;
  assign T1532 = io_invalidate ? 2'h0 : T1533;
  assign T1533 = T1528 ? T1538 : T1534;
  assign T1534 = T1536 ? T1535 : R1531;
  assign T1535 = R1531 + 2'h1;
  assign T1536 = T1543 & T1537;
  assign T1537 = R1531 < 2'h2;
  assign T1538 = R1531 - 2'h1;
  assign T1539 = io_ras_update_valid & T1540;
  assign T1540 = T1542 & T1541;
  assign T1541 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T1542 = io_ras_update_bits_isCall ^ 1'h1;
  assign T1543 = io_ras_update_valid & io_ras_update_bits_isCall;
  assign T1545 = T1546 ? io_ras_update_bits_returnAddr : R1544;
  assign T1546 = T1543 & T1547;
  assign T1547 = T1521[1'h1:1'h1];
  assign T1548 = R1524;
  assign T1549 = T1564 & T1550;
  assign T1550 = T1551 != 62'h0;
  assign T1551 = hits & useRAS;
  assign T1716 = T1552[6'h3d:1'h0];
  assign T1552 = R7 ? T1553 : T1717;
  assign T1717 = {2'h0, useRAS};
  assign T1553 = T1562 | T1554;
  assign T1554 = T1719 & T1555;
  assign T1555 = T1557 | T1718;
  assign T1718 = {2'h0, T1556};
  assign T1556 = useRAS ^ useRAS;
  assign T1557 = 1'h1 << T41;
  assign T1719 = T1558 ? 64'hffffffffffffffff : 64'h0;
  assign T1558 = T1559;
  assign T1559 = R1560;
  assign T1561 = io_btb_update_valid ? io_btb_update_bits_isReturn : R1560;
  assign T1562 = T1720 & T1563;
  assign T1563 = ~ T1555;
  assign T1720 = {2'h0, useRAS};
  assign T1564 = T1565 ^ 1'h1;
  assign T1565 = R1531 == 2'h0;
  assign T1566 = T1543 & T1550;
  assign io_resp_bits_bridx = T1567;
  assign T1567 = brIdx[io_resp_bits_entry];
  assign T1569 = R7 & T1570;
  assign T1570 = T41 < 6'h3e;
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_taken = T1571;
  assign T1571 = T1572 ? 1'h0 : io_resp_valid;
  assign T1572 = T1576 & T1573;
  assign T1573 = T1574 ^ 1'h1;
  assign T1574 = T1575 != 62'h0;
  assign T1575 = hits & isJump;
  assign T1576 = T1577 ^ 1'h1;
  assign T1577 = T8[1'h0:1'h0];
  assign io_resp_valid = T1578;
  assign T1578 = hits != 62'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
// synthesis translate_on
`endif
    if(io_btb_update_valid) begin
      R4 <= io_btb_update_bits_target;
    end
    if(reset) begin
      R7 <= 1'h0;
    end else begin
      R7 <= io_btb_update_valid;
    end
    if (T21)
      T10[T22] <= T12;
    if(T1051) begin
      R25 <= T1049;
    end else if(T31) begin
      R25 <= T28;
    end
    isJump <= T1580;
    if(reset) begin
      R42 <= 6'h0;
    end else if(T47) begin
      R42 <= T44;
    end
    if(io_btb_update_valid) begin
      R49 <= io_btb_update_bits_prediction_bits_entry;
    end
    if(io_btb_update_valid) begin
      updateHit <= io_btb_update_bits_prediction_valid;
    end
    if(io_btb_update_valid) begin
      R54 <= io_btb_update_bits_isJump;
    end
    pageValid <= T1586;
    if(reset) begin
      R75 <= 3'h0;
    end else if(T80) begin
      R75 <= T77;
    end
    if(io_btb_update_valid) begin
      R87 <= io_btb_update_bits_pc;
    end
    if (T96)
      pages[3'h5] <= T91;
    if (T101)
      pages[3'h3] <= T91;
    if (T105)
      pages[3'h1] <= T91;
    if (T112)
      pages[3'h4] <= T109;
    if (T117)
      pages[3'h2] <= T109;
    if (T121)
      pages[3'h0] <= T109;
    if (T165)
      idxPages[T41] <= T1595;
    if (T478)
      idxs[T41] <= T1606;
    idxValid <= T1607;
    if (T676)
      tgtPages[T41] <= T1611;
    if (T1062)
      tgts[T41] <= T1713;
    if(T1519) begin
      R1517 <= io_ras_update_bits_returnAddr;
    end
    if(reset) begin
      R1524 <= 1'h0;
    end else if(T1528) begin
      R1524 <= T1527;
    end else if(T1543) begin
      R1524 <= T1523;
    end
    if(reset) begin
      R1531 <= 2'h0;
    end else if(io_invalidate) begin
      R1531 <= 2'h0;
    end else if(T1528) begin
      R1531 <= T1538;
    end else if(T1536) begin
      R1531 <= T1535;
    end
    if(T1546) begin
      R1544 <= io_ras_update_bits_returnAddr;
    end
    useRAS <= T1716;
    if(io_btb_update_valid) begin
      R1560 <= io_btb_update_bits_isReturn;
    end
    if (T1569)
      brIdx[T41] <= 1'h0;
  end
endmodule

module FlowThroughSerializer(
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [135:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [3:0] io_in_bits_payload_manager_xact_id,
    input  io_in_bits_payload_uncached,
    input [1:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[135:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output io_cnt,
    output io_done
);

  wire T1;
  wire[-1:0] T0;


  assign io_done = 1'h1;
  assign io_cnt = T1;
  assign T1 = {1'h0, T0};
  assign T0 = {0{$random}};
  assign io_out_bits_payload_g_type = io_in_bits_payload_g_type;
  assign io_out_bits_payload_uncached = io_in_bits_payload_uncached;
  assign io_out_bits_payload_manager_xact_id = io_in_bits_payload_manager_xact_id;
  assign io_out_bits_payload_client_xact_id = io_in_bits_payload_client_xact_id;
  assign io_out_bits_payload_data = io_in_bits_payload_data;
  assign io_out_bits_header_dst = io_in_bits_header_dst;
  assign io_out_bits_header_src = io_in_bits_header_src;
  assign io_out_valid = io_in_valid;
  assign io_in_ready = io_out_ready;
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output io_count
);

  wire T13;
  wire[1:0] T0;
  reg  full;
  wire T14;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[3:0] T3;
  wire[7:0] T4;
  reg [7:0] ram [0:0];
  wire[7:0] T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[5:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire empty;
  wire T12;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T13;
  assign T13 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T14 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_manager_xact_id = T3;
  assign T3 = T4[2'h3:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_manager_xact_id};
  assign io_deq_bits_header_dst = T9;
  assign T9 = T4[3'h5:3'h4];
  assign io_deq_bits_header_src = T10;
  assign T10 = T4[3'h7:3'h6];
  assign io_deq_valid = T11;
  assign T11 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [12:0] io_req_bits_idx,
    input [18:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[135:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[128:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire refill_done;
  wire refill_wrap;
  wire T3;
  reg [1:0] refill_cnt;
  wire[1:0] T216;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [1:0] state;
  wire[1:0] T217;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire s2_miss;
  wire T13;
  wire s2_any_tag_hit;
  wire T14;
  wire T15;
  wire T16;
  wire s2_disparity_1;
  wire T17;
  reg  R18;
  wire T19;
  wire T20;
  wire T21;
  wire stall;
  wire T22;
  wire rdy;
  wire T23;
  wire T24;
  wire T25;
  reg  s1_valid;
  wire T218;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg  R31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  wire[6:0] T41;
  reg [12:0] s1_pgoff;
  wire[12:0] T42;
  wire T43;
  wire T44;
  reg [255:0] vb_array;
  wire[255:0] T219;
  wire[255:0] T45;
  wire[255:0] T46;
  wire[255:0] T47;
  wire[255:0] T48;
  wire[255:0] T49;
  wire[255:0] T50;
  wire[255:0] T51;
  wire[7:0] T52;
  wire[6:0] s2_idx;
  reg [31:0] s2_addr;
  wire[31:0] T53;
  wire[31:0] s1_addr;
  wire[31:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire repl_way;
  reg [15:0] R58;
  wire[15:0] T220;
  wire[15:0] T59;
  wire[15:0] T60;
  wire[14:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire[255:0] T221;
  wire T69;
  wire[255:0] T70;
  wire[255:0] T71;
  wire T72;
  wire T73;
  reg  invalidated;
  wire T74;
  wire T75;
  wire[255:0] T76;
  wire[255:0] T77;
  wire[255:0] T78;
  wire[7:0] T79;
  wire[255:0] T222;
  wire T80;
  wire[255:0] T81;
  wire[255:0] T82;
  wire T83;
  wire[255:0] T84;
  wire[255:0] T85;
  wire[255:0] T86;
  wire[7:0] T87;
  wire[255:0] T223;
  wire T88;
  wire[255:0] T89;
  wire[255:0] T90;
  wire T91;
  wire T92;
  wire s2_disparity_0;
  wire T93;
  reg  R94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg  R99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[6:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire s2_tag_hit_1;
  wire T113;
  reg  R114;
  wire T115;
  wire s1_tag_match_1;
  wire T116;
  wire[18:0] s1_tag;
  wire[18:0] T117;
  wire[18:0] T118;
  wire[37:0] T119;
  wire T133;
  wire s0_valid;
  wire T134;
  wire T135;
  wire[6:0] T131;
  wire[12:0] s0_pgoff;
  wire T132;
  wire[37:0] T120;
  wire[37:0] T121;
  wire[37:0] T122;
  wire[18:0] T123;
  wire[18:0] T224;
  wire T124;
  wire[1:0] T125;
  wire[18:0] T126;
  wire[18:0] T225;
  wire T127;
  wire[37:0] T128;
  wire[18:0] T129;
  wire[18:0] s2_tag;
  reg [6:0] tag_raddr;
  wire[6:0] T130;
  wire s2_tag_hit_0;
  wire T136;
  reg  R137;
  wire T138;
  wire s1_tag_match_0;
  wire T139;
  wire[18:0] T140;
  wire[18:0] T141;
  reg  s2_valid;
  wire T226;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire[128:0] T155;
  wire[1:0] T156;
  wire T157;
  wire[135:0] T158;
  wire[1:0] T159;
  wire[25:0] T160;
  wire[25:0] T161;
  wire T162;
  wire T163;
  wire[127:0] T164;
  wire[127:0] T165;
  reg [127:0] s2_dout_1;
  wire[127:0] T166;
  wire[127:0] T167;
  wire T180;
  wire T181;
  wire T174;
  wire T175;
  wire[8:0] T179;
  wire[127:0] T169;
  wire[127:0] T170;
  wire[127:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[8:0] T176;
  reg [8:0] R177;
  wire[8:0] T178;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[127:0] T186;
  reg [127:0] s2_dout_0;
  wire[127:0] T187;
  wire[127:0] T188;
  wire T201;
  wire T202;
  wire T195;
  wire T196;
  wire[8:0] T200;
  wire[127:0] T190;
  wire[127:0] T191;
  wire[127:0] T192;
  wire[63:0] T193;
  wire[63:0] T194;
  wire[8:0] T197;
  reg [8:0] R198;
  wire[8:0] T199;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire[31:0] T207;
  wire[31:0] T208;
  wire[31:0] s2_dout_word_1;
  wire[127:0] T209;
  wire[6:0] T210;
  wire[1:0] T211;
  wire[5:0] s2_offset;
  wire[31:0] T212;
  wire[31:0] s2_dout_word_0;
  wire[127:0] T213;
  wire[6:0] T214;
  wire[1:0] T215;
  wire s2_hit;
  wire ser_io_in_ready;
  wire ser_io_out_valid;
  wire[1:0] ser_io_out_bits_header_src;
  wire[135:0] ser_io_out_bits_payload_data;
  wire[3:0] ser_io_out_bits_payload_manager_xact_id;
  wire ser_io_out_bits_payload_uncached;
  wire[1:0] ser_io_out_bits_payload_g_type;
  wire ack_q_io_enq_ready;
  wire ack_q_io_deq_valid;
  wire[1:0] ack_q_io_deq_bits_header_src;
  wire[1:0] ack_q_io_deq_bits_header_dst;
  wire[3:0] ack_q_io_deq_bits_payload_manager_xact_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    refill_cnt = {1{$random}};
    state = {1{$random}};
    R18 = {1{$random}};
    s1_valid = {1{$random}};
    R31 = {1{$random}};
    s1_pgoff = {1{$random}};
    vb_array = {8{$random}};
    s2_addr = {1{$random}};
    R58 = {1{$random}};
    invalidated = {1{$random}};
    R94 = {1{$random}};
    R99 = {1{$random}};
    R114 = {1{$random}};
    tag_raddr = {1{$random}};
    R137 = {1{$random}};
    s2_valid = {1{$random}};
    s2_dout_1 = {4{$random}};
    R177 = {1{$random}};
    s2_dout_0 = {4{$random}};
    R198 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = refill_done & T1;
  assign T1 = ser_io_out_bits_payload_uncached | T2;
  assign T2 = ser_io_out_bits_payload_g_type != 2'h0;
  assign refill_done = T7 & refill_wrap;
  assign refill_wrap = T6 & T3;
  assign T3 = refill_cnt == 2'h3;
  assign T216 = reset ? 2'h0 : T4;
  assign T4 = T6 ? T5 : refill_cnt;
  assign T5 = refill_cnt + 2'h1;
  assign T6 = 1'h1 & ser_io_out_valid;
  assign T7 = state == 2'h3;
  assign T217 = reset ? 2'h0 : T8;
  assign T8 = T153 ? 2'h0 : T9;
  assign T9 = T151 ? 2'h3 : T10;
  assign T10 = T148 ? 2'h2 : T11;
  assign T11 = T12 ? 2'h1 : state;
  assign T12 = T147 & s2_miss;
  assign s2_miss = s2_valid & T13;
  assign T13 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T14;
  assign T14 = T112 & T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = s2_disparity_0 | s2_disparity_1;
  assign s2_disparity_1 = T17;
  assign T17 = R31 & R18;
  assign T19 = T20 ? 1'h0 : R18;
  assign T20 = T22 & T21;
  assign T21 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T22 = s1_valid & rdy;
  assign rdy = T23;
  assign T23 = T25 & T24;
  assign T24 = s2_miss ^ 1'h1;
  assign T25 = state == 2'h0;
  assign T218 = reset ? 1'h0 : T26;
  assign T26 = T30 | T27;
  assign T27 = T29 & T28;
  assign T28 = io_req_bits_kill ^ 1'h1;
  assign T29 = s1_valid & stall;
  assign T30 = io_req_valid & rdy;
  assign T32 = T20 ? T33 : R31;
  assign T33 = T92 & T34;
  assign T34 = T35;
  assign T35 = T44 & T36;
  assign T36 = T37 - 1'h1;
  assign T37 = 1'h1 << T38;
  assign T38 = T39 + 8'h1;
  assign T39 = T40 - T40;
  assign T40 = {1'h1, T41};
  assign T41 = s1_pgoff[4'hc:3'h6];
  assign T42 = T43 ? io_req_bits_idx : s1_pgoff;
  assign T43 = io_req_valid & rdy;
  assign T44 = vb_array >> T40;
  assign T219 = reset ? 256'h0 : T45;
  assign T45 = T91 ? T84 : T46;
  assign T46 = T83 ? T76 : T47;
  assign T47 = io_invalidate ? 256'h0 : T48;
  assign T48 = T72 ? T49 : vb_array;
  assign T49 = T70 | T50;
  assign T50 = T221 & T51;
  assign T51 = 1'h1 << T52;
  assign T52 = {repl_way, s2_idx};
  assign s2_idx = s2_addr[4'hc:3'h6];
  assign T53 = T55 ? s1_addr : s2_addr;
  assign s1_addr = T54;
  assign T54 = {io_req_bits_ppn, s1_pgoff};
  assign T55 = T57 & T56;
  assign T56 = stall ^ 1'h1;
  assign T57 = s1_valid & rdy;
  assign repl_way = R58[1'h0:1'h0];
  assign T220 = reset ? 16'h1 : T59;
  assign T59 = s2_miss ? T60 : R58;
  assign T60 = {T62, T61};
  assign T61 = R58[4'hf:1'h1];
  assign T62 = T64 ^ T63;
  assign T63 = R58[3'h5:3'h5];
  assign T64 = T66 ^ T65;
  assign T65 = R58[2'h3:2'h3];
  assign T66 = T68 ^ T67;
  assign T67 = R58[2'h2:2'h2];
  assign T68 = R58[1'h0:1'h0];
  assign T221 = T69 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T69 = 1'h1;
  assign T70 = vb_array & T71;
  assign T71 = ~ T51;
  assign T72 = refill_done & T73;
  assign T73 = invalidated ^ 1'h1;
  assign T74 = T147 ? 1'h0 : T75;
  assign T75 = io_invalidate ? 1'h1 : invalidated;
  assign T76 = T81 | T77;
  assign T77 = T222 & T78;
  assign T78 = 1'h1 << T79;
  assign T79 = {1'h0, s2_idx};
  assign T222 = T80 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T80 = 1'h0;
  assign T81 = vb_array & T82;
  assign T82 = ~ T78;
  assign T83 = s2_valid & s2_disparity_0;
  assign T84 = T89 | T85;
  assign T85 = T223 & T86;
  assign T86 = 1'h1 << T87;
  assign T87 = {1'h1, s2_idx};
  assign T223 = T88 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0;
  assign T88 = 1'h0;
  assign T89 = vb_array & T90;
  assign T90 = ~ T86;
  assign T91 = s2_valid & s2_disparity_1;
  assign T92 = io_invalidate ^ 1'h1;
  assign s2_disparity_0 = T93;
  assign T93 = R99 & R94;
  assign T95 = T96 ? 1'h0 : R94;
  assign T96 = T98 & T97;
  assign T97 = stall ^ 1'h1;
  assign T98 = s1_valid & rdy;
  assign T100 = T96 ? T101 : R99;
  assign T101 = T111 & T102;
  assign T102 = T103;
  assign T103 = T110 & T104;
  assign T104 = T105 - 1'h1;
  assign T105 = 1'h1 << T106;
  assign T106 = T107 + 8'h1;
  assign T107 = T108 - T108;
  assign T108 = {1'h0, T109};
  assign T109 = s1_pgoff[4'hc:3'h6];
  assign T110 = vb_array >> T108;
  assign T111 = io_invalidate ^ 1'h1;
  assign T112 = s2_tag_hit_0 | s2_tag_hit_1;
  assign s2_tag_hit_1 = T113;
  assign T113 = R31 & R114;
  assign T115 = T20 ? s1_tag_match_1 : R114;
  assign s1_tag_match_1 = T116;
  assign T116 = T117 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hd];
  assign T117 = T118[5'h12:1'h0];
  assign T118 = T119[6'h25:5'h13];
  assign T133 = T135 & s0_valid;
  assign s0_valid = io_req_valid | T134;
  assign T134 = s1_valid & stall;
  assign T135 = refill_done ^ 1'h1;
  assign T131 = s0_pgoff[4'hc:3'h6];
  assign s0_pgoff = T132 ? s1_pgoff : io_req_bits_idx;
  assign T132 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(refill_done ? s2_idx : T131),
    .RW0E(T133 || refill_done),
    .RW0W(refill_done),
    .RW0I(T128),
    .RW0M(T121),
    .RW0O(T119)
  );
  assign T121 = T122;
  assign T122 = {T126, T123};
  assign T123 = 19'h0 - T224;
  assign T224 = {18'h0, T124};
  assign T124 = T125[1'h0:1'h0];
  assign T125 = 1'h1 << repl_way;
  assign T126 = 19'h0 - T225;
  assign T225 = {18'h0, T127};
  assign T127 = T125[1'h1:1'h1];
  assign T128 = {T129, T129};
  assign T129 = s2_tag;
  assign s2_tag = s2_addr[5'h1f:4'hd];
  assign T130 = T133 ? T131 : tag_raddr;
  assign s2_tag_hit_0 = T136;
  assign T136 = R99 & R137;
  assign T138 = T96 ? s1_tag_match_0 : R137;
  assign s1_tag_match_0 = T139;
  assign T139 = T140 == s1_tag;
  assign T140 = T141[5'h12:1'h0];
  assign T141 = T119[5'h12:1'h0];
  assign T226 = reset ? 1'h0 : T142;
  assign T142 = T144 | T143;
  assign T143 = io_resp_valid & stall;
  assign T144 = T146 & T145;
  assign T145 = io_req_bits_kill ^ 1'h1;
  assign T146 = s1_valid & rdy;
  assign T147 = 2'h0 == state;
  assign T148 = T150 & T149;
  assign T149 = io_mem_acquire_ready & ack_q_io_enq_ready;
  assign T150 = 2'h1 == state;
  assign T151 = T152 & io_mem_grant_valid;
  assign T152 = 2'h2 == state;
  assign T153 = T154 & refill_done;
  assign T154 = 2'h3 == state;
  assign io_mem_finish_bits_payload_manager_xact_id = ack_q_io_deq_bits_payload_manager_xact_id;
  assign io_mem_finish_bits_header_dst = ack_q_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ack_q_io_deq_bits_header_src;
  assign io_mem_finish_valid = ack_q_io_deq_valid;
  assign io_mem_grant_ready = ser_io_in_ready;
  assign io_mem_acquire_bits_payload_subblock = T155;
  assign T155 = 129'hf;
  assign io_mem_acquire_bits_payload_a_type = T156;
  assign T156 = 2'h0;
  assign io_mem_acquire_bits_payload_uncached = T157;
  assign T157 = 1'h1;
  assign io_mem_acquire_bits_payload_data = T158;
  assign T158 = 136'h0;
  assign io_mem_acquire_bits_payload_client_xact_id = T159;
  assign T159 = 2'h0;
  assign io_mem_acquire_bits_payload_addr = T160;
  assign T160 = T161;
  assign T161 = s2_addr >> 3'h6;
//  assign io_mem_acquire_bits_header_dst = {1{$random}};
//  assign io_mem_acquire_bits_header_src = {1{$random}};
  assign io_mem_acquire_valid = T162;
  assign T162 = T163 & ack_q_io_enq_ready;
  assign T163 = state == 2'h1;
  assign io_resp_bits_datablock = T164;
  assign T164 = T186 | T165;
  assign T165 = s2_tag_hit_1 ? s2_dout_1 : 128'h0;
  assign T166 = T182 ? T167 : s2_dout_1;
  assign T180 = T181 & s0_valid;
  assign T181 = T174 ^ 1'h1;
  assign T174 = ser_io_out_valid & T175;
  assign T175 = repl_way == 1'h1;
  assign T179 = s0_pgoff[4'hc:3'h4];
  ICache_T168 T168 (
    .CLK(clk),
    .RW0A(T174 ? T176 : T179),
    .RW0E(T180 || T174),
    .RW0W(T174),
    .RW0I(T170),
    .RW0O(T167)
  );
  assign T170 = T171;
  assign T171 = {T173, T172};
  assign T172 = ser_io_out_bits_payload_data[6'h3f:1'h0];
  assign T173 = ser_io_out_bits_payload_data[8'h83:7'h44];
  assign T176 = {s2_idx, refill_cnt};
  assign T178 = T180 ? T179 : R177;
  assign T182 = T183 & s1_tag_match_1;
  assign T183 = T185 & T184;
  assign T184 = stall ^ 1'h1;
  assign T185 = s1_valid & rdy;
  assign T186 = s2_tag_hit_0 ? s2_dout_0 : 128'h0;
  assign T187 = T203 ? T188 : s2_dout_0;
  assign T201 = T202 & s0_valid;
  assign T202 = T195 ^ 1'h1;
  assign T195 = ser_io_out_valid & T196;
  assign T196 = repl_way == 1'h0;
  assign T200 = s0_pgoff[4'hc:3'h4];
  ICache_T168 T189 (
    .CLK(clk),
    .RW0A(T195 ? T197 : T200),
    .RW0E(T201 || T195),
    .RW0W(T195),
    .RW0I(T191),
    .RW0O(T188)
  );
  assign T191 = T192;
  assign T192 = {T194, T193};
  assign T193 = ser_io_out_bits_payload_data[6'h3f:1'h0];
  assign T194 = ser_io_out_bits_payload_data[8'h83:7'h44];
  assign T197 = {s2_idx, refill_cnt};
  assign T199 = T201 ? T200 : R198;
  assign T203 = T204 & s1_tag_match_0;
  assign T204 = T206 & T205;
  assign T205 = stall ^ 1'h1;
  assign T206 = s1_valid & rdy;
  assign io_resp_bits_data = T207;
  assign T207 = T212 | T208;
  assign T208 = s2_tag_hit_1 ? s2_dout_word_1 : 32'h0;
  assign s2_dout_word_1 = T209[5'h1f:1'h0];
  assign T209 = s2_dout_1 >> T210;
  assign T210 = T211 << 3'h5;
  assign T211 = s2_offset[2'h3:2'h2];
  assign s2_offset = s2_addr[3'h5:1'h0];
  assign T212 = s2_tag_hit_0 ? s2_dout_word_0 : 32'h0;
  assign s2_dout_word_0 = T213[5'h1f:1'h0];
  assign T213 = s2_dout_0 >> T214;
  assign T214 = T215 << 3'h5;
  assign T215 = s2_offset[2'h3:2'h2];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer ser(
       .io_in_ready( ser_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_in_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( ser_io_out_valid ),
       .io_out_bits_header_src( ser_io_out_bits_header_src ),
       //.io_out_bits_header_dst(  )
       .io_out_bits_payload_data( ser_io_out_bits_payload_data ),
       //.io_out_bits_payload_client_xact_id(  )
       .io_out_bits_payload_manager_xact_id( ser_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( ser_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( ser_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Queue_8 ack_q(.clk(clk), .reset(reset),
       .io_enq_ready( ack_q_io_enq_ready ),
       .io_enq_valid( T0 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( ser_io_out_bits_header_src ),
       .io_enq_bits_payload_manager_xact_id( ser_io_out_bits_payload_manager_xact_id ),
       .io_deq_ready( io_mem_finish_ready ),
       .io_deq_valid( ack_q_io_deq_valid ),
       .io_deq_bits_header_src( ack_q_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ack_q_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( ack_q_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ack_q.io_enq_bits_header_src = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T6) begin
      refill_cnt <= T5;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T153) begin
      state <= 2'h0;
    end else if(T151) begin
      state <= 2'h3;
    end else if(T148) begin
      state <= 2'h2;
    end else if(T12) begin
      state <= 2'h1;
    end
    if(T20) begin
      R18 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T26;
    end
    if(T20) begin
      R31 <= T33;
    end
    if(T43) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else if(T91) begin
      vb_array <= T84;
    end else if(T83) begin
      vb_array <= T76;
    end else if(io_invalidate) begin
      vb_array <= 256'h0;
    end else if(T72) begin
      vb_array <= T49;
    end
    if(T55) begin
      s2_addr <= s1_addr;
    end
    if(reset) begin
      R58 <= 16'h1;
    end else if(s2_miss) begin
      R58 <= T60;
    end
    if(T147) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(T96) begin
      R94 <= 1'h0;
    end
    if(T96) begin
      R99 <= T101;
    end
    if(T20) begin
      R114 <= s1_tag_match_1;
    end
    if(T133) begin
      tag_raddr <= T131;
    end
    if(T96) begin
      R137 <= s1_tag_match_0;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T142;
    end
    if(T182) begin
      s2_dout_1 <= T167;
    end
    if(T180) begin
      R177 <= T179;
    end
    if(T203) begin
      s2_dout_0 <= T188;
    end
    if(T201) begin
      R198 <= T200;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input  io_clear_hit,
    input [36:0] io_tag,
    output io_hit,
    output[7:0] io_hits,
    output[7:0] io_valid_bits,
    input  io_write,
    input [36:0] io_write_tag,
    input [2:0] io_write_addr
);

  reg [7:0] vb_array;
  wire[7:0] T47;
  wire[7:0] T0;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[7:0] T4;
  wire[7:0] T5;
  wire[7:0] T48;
  wire T6;
  wire[7:0] T7;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire T11;
  wire T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[3:0] T15;
  wire[1:0] T16;
  wire hits_0;
  wire T17;
  wire[36:0] T18;
  reg [36:0] cam_tags [7:0];
  wire[36:0] T19;
  wire T20;
  wire hits_1;
  wire T21;
  wire[36:0] T22;
  wire T23;
  wire[1:0] T24;
  wire hits_2;
  wire T25;
  wire[36:0] T26;
  wire T27;
  wire hits_3;
  wire T28;
  wire[36:0] T29;
  wire T30;
  wire[3:0] T31;
  wire[1:0] T32;
  wire hits_4;
  wire T33;
  wire[36:0] T34;
  wire T35;
  wire hits_5;
  wire T36;
  wire[36:0] T37;
  wire T38;
  wire[1:0] T39;
  wire hits_6;
  wire T40;
  wire[36:0] T41;
  wire T42;
  wire hits_7;
  wire T43;
  wire[36:0] T44;
  wire T45;
  wire T46;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_valid_bits = vb_array;
  assign T47 = reset ? 8'h0 : T0;
  assign T0 = T11 ? T9 : T1;
  assign T1 = io_clear ? 8'h0 : T2;
  assign T2 = io_write ? T3 : vb_array;
  assign T3 = T7 | T4;
  assign T4 = T48 & T5;
  assign T5 = 1'h1 << io_write_addr;
  assign T48 = T6 ? 8'hff : 8'h0;
  assign T6 = 1'h1;
  assign T7 = vb_array & T8;
  assign T8 = ~ T5;
  assign T9 = vb_array & T10;
  assign T10 = ~ io_hits;
  assign T11 = T12 & io_clear_hit;
  assign T12 = io_clear ^ 1'h1;
  assign io_hits = T13;
  assign T13 = T14;
  assign T14 = {T31, T15};
  assign T15 = {T24, T16};
  assign T16 = {hits_1, hits_0};
  assign hits_0 = T20 & T17;
  assign T17 = T18 == io_tag;
  assign T18 = cam_tags[3'h0];
  assign T20 = vb_array[1'h0:1'h0];
  assign hits_1 = T23 & T21;
  assign T21 = T22 == io_tag;
  assign T22 = cam_tags[3'h1];
  assign T23 = vb_array[1'h1:1'h1];
  assign T24 = {hits_3, hits_2};
  assign hits_2 = T27 & T25;
  assign T25 = T26 == io_tag;
  assign T26 = cam_tags[3'h2];
  assign T27 = vb_array[2'h2:2'h2];
  assign hits_3 = T30 & T28;
  assign T28 = T29 == io_tag;
  assign T29 = cam_tags[3'h3];
  assign T30 = vb_array[2'h3:2'h3];
  assign T31 = {T39, T32};
  assign T32 = {hits_5, hits_4};
  assign hits_4 = T35 & T33;
  assign T33 = T34 == io_tag;
  assign T34 = cam_tags[3'h4];
  assign T35 = vb_array[3'h4:3'h4];
  assign hits_5 = T38 & T36;
  assign T36 = T37 == io_tag;
  assign T37 = cam_tags[3'h5];
  assign T38 = vb_array[3'h5:3'h5];
  assign T39 = {hits_7, hits_6};
  assign hits_6 = T42 & T40;
  assign T40 = T41 == io_tag;
  assign T41 = cam_tags[3'h6];
  assign T42 = vb_array[3'h6:3'h6];
  assign hits_7 = T45 & T43;
  assign T43 = T44 == io_tag;
  assign T44 = cam_tags[3'h7];
  assign T45 = vb_array[3'h7:3'h7];
  assign io_hit = T46;
  assign T46 = io_hits != 8'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 8'h0;
    end else if(T11) begin
      vb_array <= T9;
    end else if(io_clear) begin
      vb_array <= 8'h0;
    end else if(io_write) begin
      vb_array <= T3;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [30:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    output io_resp_miss,
    output[7:0] io_resp_hit_idx,
    output[18:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[29:0] io_ptw_req_bits,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [18:0] io_ptw_resp_bits_ppn,
    input [5:0] io_ptw_resp_bits_perm,
    input [7:0] io_ptw_status_ip,
    input [7:0] io_ptw_status_im,
    input [6:0] io_ptw_status_zero,
    input  io_ptw_status_er,
    input  io_ptw_status_vm,
    input  io_ptw_status_s64,
    input  io_ptw_status_u64,
    input  io_ptw_status_ef,
    input  io_ptw_status_pei,
    input  io_ptw_status_ei,
    input  io_ptw_status_ps,
    input  io_ptw_status_s,
    input  io_ptw_invalidate,
    input  io_ptw_sret
);

  reg [2:0] r_refill_waddr;
  wire[2:0] T0;
  wire[2:0] repl_waddr;
  wire[2:0] T1;
  wire[3:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  reg [7:0] R9;
  wire[7:0] T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[7:0] T13;
  wire[14:0] T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T184;
  wire[1:0] T185;
  wire T186;
  wire[1:0] T187;
  wire[1:0] T188;
  wire[3:0] T189;
  wire[3:0] T190;
  wire[3:0] T191;
  wire[1:0] T192;
  wire T193;
  wire T194;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[10:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire tlb_hit;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire[1:0] T40;
  wire T41;
  wire[2:0] T195;
  wire[2:0] T196;
  wire[2:0] T197;
  wire[2:0] T198;
  wire[2:0] T199;
  wire[2:0] T200;
  wire[2:0] T201;
  wire T202;
  wire[7:0] T42;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire has_invalid_entry;
  wire T43;
  wire T44;
  wire tlb_miss;
  wire T45;
  wire bad_va;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[36:0] T209;
  reg [37:0] r_refill_tag;
  wire[37:0] T51;
  wire[37:0] lookup_tag;
  wire[37:0] T52;
  wire T53;
  wire T54;
  reg [1:0] state;
  wire[1:0] T210;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[36:0] T211;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[29:0] T212;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[7:0] T77;
  reg [7:0] ux_array;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T213;
  wire T82;
  wire T83;
  wire[5:0] T84;
  wire[5:0] T214;
  wire T85;
  wire T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire T89;
  wire[7:0] T90;
  reg [7:0] sx_array;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire[7:0] T215;
  wire T95;
  wire T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[7:0] T104;
  reg [7:0] uw_array;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[7:0] T216;
  wire T109;
  wire T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire T113;
  wire[7:0] T114;
  reg [7:0] sw_array;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T217;
  wire T119;
  wire T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire[7:0] T128;
  reg [7:0] ur_array;
  wire[7:0] T129;
  wire[7:0] T130;
  wire[7:0] T131;
  wire[7:0] T132;
  wire[7:0] T218;
  wire T133;
  wire T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire T137;
  wire[7:0] T138;
  reg [7:0] sr_array;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[7:0] T141;
  wire[7:0] T142;
  wire[7:0] T219;
  wire T143;
  wire T144;
  wire[7:0] T145;
  wire[7:0] T146;
  wire[18:0] T147;
  wire[18:0] T148;
  wire[18:0] T149;
  wire[18:0] T150;
  wire[18:0] T151;
  reg [18:0] tag_ram [7:0];
  wire[18:0] T152;
  wire T153;
  wire[18:0] T154;
  wire[18:0] T155;
  wire[18:0] T156;
  wire T157;
  wire[18:0] T158;
  wire[18:0] T159;
  wire[18:0] T160;
  wire T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[18:0] T164;
  wire T165;
  wire[18:0] T166;
  wire[18:0] T167;
  wire[18:0] T168;
  wire T169;
  wire[18:0] T170;
  wire[18:0] T171;
  wire[18:0] T172;
  wire T173;
  wire[18:0] T174;
  wire[18:0] T175;
  wire[18:0] T176;
  wire T177;
  wire[18:0] T178;
  wire[18:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire tag_cam_io_hit;
  wire[7:0] tag_cam_io_hits;
  wire[7:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R9 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    ux_array = {1{$random}};
    sx_array = {1{$random}};
    uw_array = {1{$random}};
    sw_array = {1{$random}};
    ur_array = {1{$random}};
    sr_array = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T44 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T195 : T1;
  assign T1 = T2[2'h2:1'h0];
  assign T2 = {T33, T3};
  assign T3 = T8 & T4;
  assign T4 = T5 - 1'h1;
  assign T5 = 1'h1 << T6;
  assign T6 = T7 + 3'h1;
  assign T7 = T33 - T33;
  assign T8 = R9 >> T33;
  assign T10 = T32 ? T11 : R9;
  assign T11 = T21 | T12;
  assign T12 = T20 ? 8'h0 : T13;
  assign T13 = T14[3'h7:1'h0];
  assign T14 = 8'h1 << T15;
  assign T15 = {T18, T16};
  assign T16 = T184[1'h1:1'h1];
  assign T184 = {T194, T185};
  assign T185 = {T193, T186};
  assign T186 = T187[1'h1:1'h1];
  assign T187 = T192 | T188;
  assign T188 = T189[1'h1:1'h0];
  assign T189 = T191 | T190;
  assign T190 = tag_cam_io_hits[2'h3:1'h0];
  assign T191 = tag_cam_io_hits[3'h7:3'h4];
  assign T192 = T189[2'h3:2'h2];
  assign T193 = T192 != 2'h0;
  assign T194 = T191 != 4'h0;
  assign T18 = {1'h1, T19};
  assign T19 = T184[2'h2:2'h2];
  assign T20 = T184[1'h0:1'h0];
  assign T21 = T23 & T22;
  assign T22 = ~ T13;
  assign T23 = T27 | T24;
  assign T24 = T16 ? 8'h0 : T25;
  assign T25 = T26[3'h7:1'h0];
  assign T26 = 8'h1 << T18;
  assign T27 = T29 & T28;
  assign T28 = ~ T25;
  assign T29 = T31 | T30;
  assign T30 = T19 ? 8'h0 : 8'h2;
  assign T31 = R9 & 8'hfd;
  assign T32 = io_req_valid & tlb_hit;
  assign tlb_hit = io_ptw_status_vm & tag_cam_io_hit;
  assign T33 = {T40, T34};
  assign T34 = T39 & T35;
  assign T35 = T36 - 1'h1;
  assign T36 = 1'h1 << T37;
  assign T37 = T38 + 2'h1;
  assign T38 = T40 - T40;
  assign T39 = R9 >> T40;
  assign T40 = {1'h1, T41};
  assign T41 = R9[1'h1:1'h1];
  assign T195 = T208 ? 1'h0 : T196;
  assign T196 = T207 ? 1'h1 : T197;
  assign T197 = T206 ? 2'h2 : T198;
  assign T198 = T205 ? 2'h3 : T199;
  assign T199 = T204 ? 3'h4 : T200;
  assign T200 = T203 ? 3'h5 : T201;
  assign T201 = T202 ? 3'h6 : 3'h7;
  assign T202 = T42[3'h6:3'h6];
  assign T42 = ~ tag_cam_io_valid_bits;
  assign T203 = T42[3'h5:3'h5];
  assign T204 = T42[3'h4:3'h4];
  assign T205 = T42[2'h3:2'h3];
  assign T206 = T42[2'h2:2'h2];
  assign T207 = T42[1'h1:1'h1];
  assign T208 = T42[1'h0:1'h0];
  assign has_invalid_entry = T43 ^ 1'h1;
  assign T43 = tag_cam_io_valid_bits == 8'hff;
  assign T44 = T50 & tlb_miss;
  assign tlb_miss = T48 & T45;
  assign T45 = bad_va ^ 1'h1;
  assign bad_va = T47 != T46;
  assign T46 = io_req_bits_vpn[5'h1d:5'h1d];
  assign T47 = io_req_bits_vpn[5'h1e:5'h1e];
  assign T48 = io_ptw_status_vm & T49;
  assign T49 = tag_cam_io_hit ^ 1'h1;
  assign T50 = io_req_ready & io_req_valid;
  assign T209 = r_refill_tag[6'h24:1'h0];
  assign T51 = T44 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T52;
  assign T52 = {io_req_bits_asid, io_req_bits_vpn};
  assign T53 = T54 & io_ptw_resp_valid;
  assign T54 = state == 2'h2;
  assign T210 = reset ? 2'h0 : T55;
  assign T55 = io_ptw_resp_valid ? 2'h0 : T56;
  assign T56 = T65 ? 2'h3 : T57;
  assign T57 = T64 ? 2'h3 : T58;
  assign T58 = T63 ? 2'h2 : T59;
  assign T59 = T61 ? 2'h0 : T60;
  assign T60 = T44 ? 2'h1 : state;
  assign T61 = T62 & io_ptw_invalidate;
  assign T62 = state == 2'h1;
  assign T63 = T62 & io_ptw_req_ready;
  assign T64 = T63 & io_ptw_invalidate;
  assign T65 = T66 & io_ptw_invalidate;
  assign T66 = state == 2'h2;
  assign T211 = lookup_tag[6'h24:1'h0];
  assign T67 = T70 & T68;
  assign T68 = io_req_bits_instruction ? io_resp_xcpt_if : T69;
  assign T69 = io_resp_xcpt_ld & io_resp_xcpt_st;
  assign T70 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits = T212;
  assign T212 = r_refill_tag[5'h1d:1'h0];
  assign io_ptw_req_valid = T71;
  assign T71 = state == 2'h1;
  assign io_resp_xcpt_if = T72;
  assign T72 = bad_va | T73;
  assign T73 = tlb_hit & T74;
  assign T74 = T75 ^ 1'h1;
  assign T75 = io_ptw_status_s ? T89 : T76;
  assign T76 = T77 != 8'h0;
  assign T77 = ux_array & tag_cam_io_hits;
  assign T78 = io_ptw_resp_valid ? T79 : ux_array;
  assign T79 = T87 | T80;
  assign T80 = T213 & T81;
  assign T81 = 1'h1 << r_refill_waddr;
  assign T213 = T82 ? 8'hff : 8'h0;
  assign T82 = T83;
  assign T83 = T84[2'h2:2'h2];
  assign T84 = T214 & io_ptw_resp_bits_perm;
  assign T214 = T85 ? 6'h3f : 6'h0;
  assign T85 = T86;
  assign T86 = io_ptw_resp_bits_error ^ 1'h1;
  assign T87 = ux_array & T88;
  assign T88 = ~ T81;
  assign T89 = T90 != 8'h0;
  assign T90 = sx_array & tag_cam_io_hits;
  assign T91 = io_ptw_resp_valid ? T92 : sx_array;
  assign T92 = T97 | T93;
  assign T93 = T215 & T94;
  assign T94 = 1'h1 << r_refill_waddr;
  assign T215 = T95 ? 8'hff : 8'h0;
  assign T95 = T96;
  assign T96 = T84[3'h5:3'h5];
  assign T97 = sx_array & T98;
  assign T98 = ~ T94;
  assign io_resp_xcpt_st = T99;
  assign T99 = bad_va | T100;
  assign T100 = tlb_hit & T101;
  assign T101 = T102 ^ 1'h1;
  assign T102 = io_ptw_status_s ? T113 : T103;
  assign T103 = T104 != 8'h0;
  assign T104 = uw_array & tag_cam_io_hits;
  assign T105 = io_ptw_resp_valid ? T106 : uw_array;
  assign T106 = T111 | T107;
  assign T107 = T216 & T108;
  assign T108 = 1'h1 << r_refill_waddr;
  assign T216 = T109 ? 8'hff : 8'h0;
  assign T109 = T110;
  assign T110 = T84[1'h1:1'h1];
  assign T111 = uw_array & T112;
  assign T112 = ~ T108;
  assign T113 = T114 != 8'h0;
  assign T114 = sw_array & tag_cam_io_hits;
  assign T115 = io_ptw_resp_valid ? T116 : sw_array;
  assign T116 = T121 | T117;
  assign T117 = T217 & T118;
  assign T118 = 1'h1 << r_refill_waddr;
  assign T217 = T119 ? 8'hff : 8'h0;
  assign T119 = T120;
  assign T120 = T84[3'h4:3'h4];
  assign T121 = sw_array & T122;
  assign T122 = ~ T118;
  assign io_resp_xcpt_ld = T123;
  assign T123 = bad_va | T124;
  assign T124 = tlb_hit & T125;
  assign T125 = T126 ^ 1'h1;
  assign T126 = io_ptw_status_s ? T137 : T127;
  assign T127 = T128 != 8'h0;
  assign T128 = ur_array & tag_cam_io_hits;
  assign T129 = io_ptw_resp_valid ? T130 : ur_array;
  assign T130 = T135 | T131;
  assign T131 = T218 & T132;
  assign T132 = 1'h1 << r_refill_waddr;
  assign T218 = T133 ? 8'hff : 8'h0;
  assign T133 = T134;
  assign T134 = T84[1'h0:1'h0];
  assign T135 = ur_array & T136;
  assign T136 = ~ T132;
  assign T137 = T138 != 8'h0;
  assign T138 = sr_array & tag_cam_io_hits;
  assign T139 = io_ptw_resp_valid ? T140 : sr_array;
  assign T140 = T145 | T141;
  assign T141 = T219 & T142;
  assign T142 = 1'h1 << r_refill_waddr;
  assign T219 = T143 ? 8'hff : 8'h0;
  assign T143 = T144;
  assign T144 = T84[2'h3:2'h3];
  assign T145 = sr_array & T146;
  assign T146 = ~ T142;
  assign io_resp_ppn = T147;
  assign T147 = T181 ? T149 : T148;
  assign T148 = io_req_bits_vpn[5'h12:1'h0];
  assign T149 = T154 | T150;
  assign T150 = T153 ? T151 : 19'h0;
  assign T151 = tag_ram[3'h7];
  assign T153 = tag_cam_io_hits[3'h7:3'h7];
  assign T154 = T158 | T155;
  assign T155 = T157 ? T156 : 19'h0;
  assign T156 = tag_ram[3'h6];
  assign T157 = tag_cam_io_hits[3'h6:3'h6];
  assign T158 = T162 | T159;
  assign T159 = T161 ? T160 : 19'h0;
  assign T160 = tag_ram[3'h5];
  assign T161 = tag_cam_io_hits[3'h5:3'h5];
  assign T162 = T166 | T163;
  assign T163 = T165 ? T164 : 19'h0;
  assign T164 = tag_ram[3'h4];
  assign T165 = tag_cam_io_hits[3'h4:3'h4];
  assign T166 = T170 | T167;
  assign T167 = T169 ? T168 : 19'h0;
  assign T168 = tag_ram[3'h3];
  assign T169 = tag_cam_io_hits[2'h3:2'h3];
  assign T170 = T174 | T171;
  assign T171 = T173 ? T172 : 19'h0;
  assign T172 = tag_ram[3'h2];
  assign T173 = tag_cam_io_hits[2'h2:2'h2];
  assign T174 = T178 | T175;
  assign T175 = T177 ? T176 : 19'h0;
  assign T176 = tag_ram[3'h1];
  assign T177 = tag_cam_io_hits[1'h1:1'h1];
  assign T178 = T180 ? T179 : 19'h0;
  assign T179 = tag_ram[3'h0];
  assign T180 = tag_cam_io_hits[1'h0:1'h0];
  assign T181 = io_ptw_status_vm & T182;
  assign T182 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T183;
  assign T183 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( io_ptw_invalidate ),
       .io_clear_hit( T67 ),
       .io_tag( T211 ),
       .io_hit( tag_cam_io_hit ),
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T53 ),
       .io_write_tag( T209 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T44) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T32) begin
      R9 <= T11;
    end
    if(T44) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T65) begin
      state <= 2'h3;
    end else if(T64) begin
      state <= 2'h3;
    end else if(T63) begin
      state <= 2'h2;
    end else if(T61) begin
      state <= 2'h0;
    end else if(T44) begin
      state <= 2'h1;
    end
    if(io_ptw_resp_valid) begin
      ux_array <= T79;
    end
    if(io_ptw_resp_valid) begin
      sx_array <= T92;
    end
    if(io_ptw_resp_valid) begin
      uw_array <= T106;
    end
    if(io_ptw_resp_valid) begin
      sw_array <= T116;
    end
    if(io_ptw_resp_valid) begin
      ur_array <= T130;
    end
    if(io_ptw_resp_valid) begin
      sr_array <= T140;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [43:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[43:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data_0,
    output io_cpu_resp_bits_mask,
    output io_cpu_resp_bits_xcpt_ma,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output io_cpu_btb_resp_bits_mask,
    output io_cpu_btb_resp_bits_bridx,
    output[42:0] io_cpu_btb_resp_bits_target,
    output[5:0] io_cpu_btb_resp_bits_entry,
    output[6:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input  io_cpu_btb_update_bits_prediction_bits_mask,
    input  io_cpu_btb_update_bits_prediction_bits_bridx,
    input [42:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_btb_update_bits_pc,
    input [42:0] io_cpu_btb_update_bits_target,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isReturn,
    input [42:0] io_cpu_btb_update_bits_br_pc,
    input  io_cpu_bht_update_valid,
    input  io_cpu_bht_update_bits_prediction_valid,
    input  io_cpu_bht_update_bits_prediction_bits_taken,
    input  io_cpu_bht_update_bits_prediction_bits_mask,
    input  io_cpu_bht_update_bits_prediction_bits_bridx,
    input [42:0] io_cpu_bht_update_bits_prediction_bits_target,
    input [5:0] io_cpu_bht_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_bht_update_bits_pc,
    input  io_cpu_bht_update_bits_taken,
    input  io_cpu_bht_update_bits_mispredict,
    input  io_cpu_ras_update_valid,
    input  io_cpu_ras_update_bits_isCall,
    input  io_cpu_ras_update_bits_isReturn,
    input [42:0] io_cpu_ras_update_bits_returnAddr,
    input  io_cpu_ras_update_bits_prediction_valid,
    input  io_cpu_ras_update_bits_prediction_bits_taken,
    input  io_cpu_ras_update_bits_prediction_bits_mask,
    input  io_cpu_ras_update_bits_prediction_bits_bridx,
    input [42:0] io_cpu_ras_update_bits_prediction_bits_target,
    input [5:0] io_cpu_ras_update_bits_prediction_bits_entry,
    input [6:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    input  io_cpu_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[135:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[128:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id
);

  wire[30:0] T0;
  wire[43:0] s1_pc;
  reg [43:0] s1_pc_;
  wire[43:0] T1;
  wire[43:0] T2;
  wire[43:0] npc;
  wire[43:0] T3;
  wire[43:0] predicted_npc;
  wire[43:0] ntpc;
  wire[42:0] T4;
  wire[40:0] T5;
  wire[43:0] ntpc_0;
  wire T6;
  wire T7;
  wire T8;
  wire[43:0] btbTarget;
  wire T9;
  reg [43:0] s2_pc;
  wire[43:0] T69;
  wire[43:0] T10;
  wire T11;
  wire T12;
  wire icmiss;
  wire T13;
  reg  s2_valid;
  wire T70;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire stall;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  reg  s1_same_block;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire s0_same_block;
  wire T28;
  wire[43:0] T29;
  wire[43:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[12:0] T71;
  wire[43:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[42:0] T72;
  wire[43:0] T45;
  wire T46;
  wire T47;
  wire T48;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T49;
  wire T50;
  reg [6:0] s2_btb_resp_bits_bht_history;
  wire[6:0] T51;
  reg [5:0] s2_btb_resp_bits_entry;
  wire[5:0] T52;
  reg [42:0] s2_btb_resp_bits_target;
  wire[42:0] T53;
  reg  s2_btb_resp_bits_bridx;
  wire T54;
  reg  s2_btb_resp_bits_mask;
  wire T55;
  reg  s2_btb_resp_bits_taken;
  wire T56;
  reg  s2_btb_resp_valid;
  wire T73;
  wire T57;
  reg  s2_xcpt_if;
  wire T74;
  wire T58;
  wire T59;
  wire[1:0] T60;
  wire T75;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T76;
  wire[31:0] T63;
  wire[127:0] fetch_data;
  wire[6:0] T64;
  wire[1:0] T65;
  wire[43:0] T66;
  wire T67;
  wire T68;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire btb_io_resp_bits_mask;
  wire btb_io_resp_bits_bridx;
  wire[42:0] btb_io_resp_bits_target;
  wire[5:0] btb_io_resp_bits_entry;
  wire[6:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[135:0] icache_io_mem_acquire_bits_payload_data;
  wire icache_io_mem_acquire_bits_payload_uncached;
  wire[1:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[128:0] icache_io_mem_acquire_bits_payload_subblock;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[3:0] icache_io_mem_finish_bits_payload_manager_xact_id;
  wire tlb_io_resp_miss;
  wire[18:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[29:0] tlb_io_ptw_req_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_bridx = {1{$random}};
    s2_btb_resp_bits_mask = {1{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = s1_pc >> 4'hd;
  assign s1_pc = s1_pc_ & 44'hffffffffffe;
  assign T1 = io_cpu_req_valid ? io_cpu_req_bits_pc : T2;
  assign T2 = T17 ? npc : s1_pc_;
  assign npc = T3;
  assign T3 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : ntpc;
  assign ntpc = {T6, T4};
  assign T4 = {T5, 2'h0};
  assign T5 = ntpc_0[6'h2a:2'h2];
  assign ntpc_0 = s1_pc + 44'h4;
  assign T6 = T8 & T7;
  assign T7 = ntpc_0[6'h2a:6'h2a];
  assign T8 = s1_pc[6'h2a:6'h2a];
  assign btbTarget = {T9, btb_io_resp_bits_target};
  assign T9 = btb_io_resp_bits_target[6'h2a:6'h2a];
  assign T69 = reset ? 44'h2000 : T10;
  assign T10 = T11 ? s1_pc : s2_pc;
  assign T11 = T17 & T12;
  assign T12 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T13;
  assign T13 = icache_io_resp_valid ^ 1'h1;
  assign T70 = reset ? 1'h1 : T14;
  assign T14 = io_cpu_req_valid ? 1'h0 : T15;
  assign T15 = T17 ? T16 : s2_valid;
  assign T16 = icmiss ^ 1'h1;
  assign T17 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T18;
  assign T18 = io_cpu_resp_ready ^ 1'h1;
  assign T19 = T21 & T20;
  assign T20 = icmiss ^ 1'h1;
  assign T21 = stall ^ 1'h1;
  assign T22 = T36 & T23;
  assign T23 = s1_same_block ^ 1'h1;
  assign T24 = io_cpu_req_valid ? 1'h0 : T25;
  assign T25 = T17 ? T26 : s1_same_block;
  assign T26 = s0_same_block & T27;
  assign T27 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T31 & T28;
  assign T28 = T30 == T29;
  assign T29 = s1_pc & 44'h10;
  assign T30 = ntpc & 44'h10;
  assign T31 = T33 & T32;
  assign T32 = btb_io_resp_bits_taken ^ 1'h1;
  assign T33 = T35 & T34;
  assign T34 = io_cpu_req_valid ^ 1'h1;
  assign T35 = icmiss ^ 1'h1;
  assign T36 = stall ^ 1'h1;
  assign T37 = T38 | io_cpu_ptw_invalidate;
  assign T38 = T39 | icmiss;
  assign T39 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T71 = T40[4'hc:1'h0];
  assign T40 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T41 = T43 & T42;
  assign T42 = s0_same_block ^ 1'h1;
  assign T43 = stall ^ 1'h1;
  assign T44 = io_cpu_invalidate | io_cpu_ptw_invalidate;
  assign T72 = T45[6'h2a:1'h0];
  assign T45 = s1_pc & 44'hffffffffffc;
  assign T46 = T48 & T47;
  assign T47 = icmiss ^ 1'h1;
  assign T48 = stall ^ 1'h1;
  assign io_mem_finish_bits_payload_manager_xact_id = icache_io_mem_finish_bits_payload_manager_xact_id;
  assign io_mem_finish_bits_header_dst = icache_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = icache_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = icache_io_mem_finish_valid;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_payload_subblock = icache_io_mem_acquire_bits_payload_subblock;
  assign io_mem_acquire_bits_payload_a_type = icache_io_mem_acquire_bits_payload_a_type;
  assign io_mem_acquire_bits_payload_uncached = icache_io_mem_acquire_bits_payload_uncached;
  assign io_mem_acquire_bits_payload_data = icache_io_mem_acquire_bits_payload_data;
  assign io_mem_acquire_bits_payload_client_xact_id = icache_io_mem_acquire_bits_payload_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = icache_io_mem_acquire_bits_payload_addr;
//  assign io_mem_acquire_bits_header_dst = {1{$random}};
//  assign io_mem_acquire_bits_header_src = {1{$random}};
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cpu_ptw_req_bits = tlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T49 = T50 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T50 = T11 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T51 = T50 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T52 = T50 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T53 = T50 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign T54 = T50 ? btb_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign T55 = T50 ? btb_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T56 = T50 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T73 = reset ? 1'h0 : T57;
  assign T57 = T11 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T74 = reset ? 1'h0 : T58;
  assign T58 = T11 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_xcpt_ma = T59;
  assign T59 = T60 != 2'h0;
  assign T60 = s2_pc[1'h1:1'h0];
  assign io_cpu_resp_bits_mask = T75;
  assign T75 = T61[1'h0:1'h0];
  assign T61 = s2_btb_resp_valid ? T62 : 2'h3;
  assign T62 = 2'h3 & T76;
  assign T76 = {1'h0, s2_btb_resp_bits_mask};
  assign io_cpu_resp_bits_data_0 = T63;
  assign T63 = fetch_data[5'h1f:1'h0];
  assign fetch_data = icache_io_resp_bits_datablock >> T64;
  assign T64 = T65 << 3'h5;
  assign T65 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = T66;
  assign T66 = s2_pc & 44'hffffffffffc;
  assign io_cpu_resp_valid = T67;
  assign T67 = s2_valid & T68;
  assign T68 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T46 ),
       .io_req_bits_addr( T72 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_mask( btb_io_resp_bits_mask ),
       .io_resp_bits_bridx( btb_io_resp_bits_bridx ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_btb_update_valid( io_cpu_btb_update_valid ),
       .io_btb_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_btb_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_btb_update_bits_prediction_bits_mask( io_cpu_btb_update_bits_prediction_bits_mask ),
       .io_btb_update_bits_prediction_bits_bridx( io_cpu_btb_update_bits_prediction_bits_bridx ),
       .io_btb_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_btb_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_btb_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_btb_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_btb_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_btb_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_btb_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_btb_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_btb_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_btb_update_bits_br_pc( io_cpu_btb_update_bits_br_pc ),
       .io_bht_update_valid( io_cpu_bht_update_valid ),
       .io_bht_update_bits_prediction_valid( io_cpu_bht_update_bits_prediction_valid ),
       .io_bht_update_bits_prediction_bits_taken( io_cpu_bht_update_bits_prediction_bits_taken ),
       .io_bht_update_bits_prediction_bits_mask( io_cpu_bht_update_bits_prediction_bits_mask ),
       .io_bht_update_bits_prediction_bits_bridx( io_cpu_bht_update_bits_prediction_bits_bridx ),
       .io_bht_update_bits_prediction_bits_target( io_cpu_bht_update_bits_prediction_bits_target ),
       .io_bht_update_bits_prediction_bits_entry( io_cpu_bht_update_bits_prediction_bits_entry ),
       .io_bht_update_bits_prediction_bits_bht_history( io_cpu_bht_update_bits_prediction_bits_bht_history ),
       .io_bht_update_bits_prediction_bits_bht_value( io_cpu_bht_update_bits_prediction_bits_bht_value ),
       .io_bht_update_bits_pc( io_cpu_bht_update_bits_pc ),
       .io_bht_update_bits_taken( io_cpu_bht_update_bits_taken ),
       .io_bht_update_bits_mispredict( io_cpu_bht_update_bits_mispredict ),
       .io_ras_update_valid( io_cpu_ras_update_valid ),
       .io_ras_update_bits_isCall( io_cpu_ras_update_bits_isCall ),
       .io_ras_update_bits_isReturn( io_cpu_ras_update_bits_isReturn ),
       .io_ras_update_bits_returnAddr( io_cpu_ras_update_bits_returnAddr ),
       .io_ras_update_bits_prediction_valid( io_cpu_ras_update_bits_prediction_valid ),
       .io_ras_update_bits_prediction_bits_taken( io_cpu_ras_update_bits_prediction_bits_taken ),
       .io_ras_update_bits_prediction_bits_mask( io_cpu_ras_update_bits_prediction_bits_mask ),
       .io_ras_update_bits_prediction_bits_bridx( io_cpu_ras_update_bits_prediction_bits_bridx ),
       .io_ras_update_bits_prediction_bits_target( io_cpu_ras_update_bits_prediction_bits_target ),
       .io_ras_update_bits_prediction_bits_entry( io_cpu_ras_update_bits_prediction_bits_entry ),
       .io_ras_update_bits_prediction_bits_bht_history( io_cpu_ras_update_bits_prediction_bits_bht_history ),
       .io_ras_update_bits_prediction_bits_bht_value( io_cpu_ras_update_bits_prediction_bits_bht_value ),
       .io_invalidate( T44 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T41 ),
       .io_req_bits_idx( T71 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T37 ),
       .io_resp_ready( T22 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( icache_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( icache_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( icache_io_mem_finish_bits_payload_manager_xact_id )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T19 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T0 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_resp_miss( tlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits( tlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T17) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 44'h2000;
    end else if(T11) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T17) begin
      s2_valid <= T16;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T17) begin
      s1_same_block <= T26;
    end
    if(T50) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T50) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T50) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T50) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T50) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if(T50) begin
      s2_btb_resp_bits_mask <= btb_io_resp_bits_mask;
    end
    if(T50) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T11) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T11) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [18:0] io_req_bits_tag,
    input [6:0] io_req_bits_idx,
    input [3:0] io_req_bits_way_en,
    input [1:0] io_req_bits_client_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output[3:0] io_data_req_bits_way_en,
    output[12:0] io_data_req_bits_addr,
    input [135:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr,
    output[1:0] io_release_bits_client_xact_id,
    output[135:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg [1:0] req_client_xact_id;
  wire[1:0] T2;
  wire[25:0] T3;
  wire[25:0] T4;
  reg [6:0] req_idx;
  wire[6:0] T5;
  reg [18:0] req_tag;
  wire[18:0] T6;
  wire T7;
  reg  r2_data_req_fired;
  wire T36;
  wire T8;
  wire T9;
  reg  r1_data_req_fired;
  wire T37;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg  active;
  wire T38;
  wire T19;
  wire T20;
  wire T21;
  reg [2:0] cnt;
  wire[2:0] T39;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T40;
  wire[1:0] T27;
  wire T28;
  wire T29;
  wire[12:0] T30;
  wire[8:0] T31;
  wire[1:0] T32;
  reg [3:0] req_way_en;
  wire[3:0] T33;
  wire fire;
  wire T34;
  wire T35;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_idx = {1{$random}};
    req_tag = {1{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    cnt = {1{$random}};
    req_way_en = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_data = io_data_resp;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T2 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr = T3;
  assign T3 = T4;
  assign T4 = {req_tag, req_idx};
  assign T5 = T1 ? io_req_bits_idx : req_idx;
  assign T6 = T1 ? io_req_bits_tag : req_tag;
  assign io_release_valid = T7;
  assign T7 = active & r2_data_req_fired;
  assign T36 = reset ? 1'h0 : T8;
  assign T8 = T17 ? 1'h0 : T9;
  assign T9 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T37 = reset ? 1'h0 : T10;
  assign T10 = T17 ? 1'h0 : T11;
  assign T11 = T13 ? 1'h1 : T12;
  assign T12 = active ? 1'h0 : r1_data_req_fired;
  assign T13 = active & T14;
  assign T14 = T16 & T15;
  assign T15 = io_meta_read_ready & io_meta_read_valid;
  assign T16 = io_data_req_ready & io_data_req_valid;
  assign T17 = T7 & T18;
  assign T18 = io_release_ready ^ 1'h1;
  assign T38 = reset ? 1'h0 : T19;
  assign T19 = T1 ? 1'h1 : T20;
  assign T20 = T28 ? T21 : active;
  assign T21 = cnt < 3'h4;
  assign T39 = reset ? 3'h0 : T22;
  assign T22 = T1 ? 3'h0 : T23;
  assign T23 = T17 ? T26 : T24;
  assign T24 = T13 ? T25 : cnt;
  assign T25 = cnt + 3'h1;
  assign T26 = cnt - T40;
  assign T40 = {1'h0, T27};
  assign T27 = r1_data_req_fired ? 2'h2 : 2'h1;
  assign T28 = T7 & T29;
  assign T29 = r1_data_req_fired ^ 1'h1;
  assign io_data_req_bits_addr = T30;
  assign T30 = T31 << 3'h4;
  assign T31 = {req_idx, T32};
  assign T32 = cnt[1'h1:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T33 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T34;
  assign T34 = cnt < 3'h4;
  assign io_meta_read_bits_tag = req_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T35;
  assign T35 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_idx <= io_req_bits_idx;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(T17) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T17) begin
      r1_data_req_fired <= 1'h0;
    end else if(T13) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T28) begin
      active <= T21;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else if(T1) begin
      cnt <= 3'h0;
    end else if(T17) begin
      cnt <= T26;
    end else if(T13) begin
      cnt <= T25;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr,
    input [1:0] io_req_bits_p_type,
    input [1:0] io_req_bits_client_xact_id,
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr,
    output[1:0] io_rep_bits_client_xact_id,
    output[135:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    input [3:0] io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_line_state_state
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  reg [1:0] req_p_type;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [3:0] state;
  wire[3:0] T91;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  reg [1:0] line_state_state;
  wire[1:0] T29;
  wire T30;
  wire hit;
  reg [3:0] way_en;
  wire[3:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  reg [1:0] req_client_xact_id;
  wire[1:0] T50;
  wire[6:0] T92;
  reg [25:0] req_addr;
  wire[25:0] T51;
  wire[18:0] T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[18:0] T61;
  wire[6:0] T93;
  wire T62;
  wire[18:0] T63;
  wire[6:0] T94;
  wire T64;
  wire[2:0] T65;
  wire[2:0] T66;
  wire[2:0] T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire[135:0] T82;
  wire[1:0] T83;
  wire[25:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_p_type = {1{$random}};
    state = {1{$random}};
    line_state_state = {1{$random}};
    way_en = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_wb_req_bits_r_type = T0;
  assign T0 = T47 ? T41 : T1;
  assign T1 = T40 ? 3'h4 : T2;
  assign T2 = T39 ? 3'h5 : T3;
  assign T3 = T4 ? 3'h6 : 3'h4;
  assign T4 = req_p_type == 2'h2;
  assign T5 = T6 ? io_req_bits_p_type : req_p_type;
  assign T6 = T7 & io_req_valid;
  assign T7 = state == 4'h1;
  assign T91 = reset ? 4'h1 : T8;
  assign T8 = T38 ? 4'h1 : T9;
  assign T9 = T6 ? 4'h2 : T10;
  assign T10 = T36 ? 4'h3 : T11;
  assign T11 = T35 ? 4'h4 : T12;
  assign T12 = T33 ? 4'h2 : T13;
  assign T13 = T32 ? 4'h5 : T14;
  assign T14 = T30 ? T27 : T15;
  assign T15 = T25 ? 4'h1 : T16;
  assign T16 = T23 ? 4'h7 : T17;
  assign T17 = T21 ? 4'h8 : T18;
  assign T18 = T19 ? 4'h1 : state;
  assign T19 = T20 & io_meta_write_ready;
  assign T20 = state == 4'h8;
  assign T21 = T22 & io_wb_req_ready;
  assign T22 = state == 4'h7;
  assign T23 = T24 & io_wb_req_ready;
  assign T24 = state == 4'h6;
  assign T25 = T26 & io_rep_ready;
  assign T26 = state == 4'h5;
  assign T27 = T28 ? 4'h6 : 4'h8;
  assign T28 = line_state_state == 2'h2;
  assign T29 = T32 ? io_line_state_state : line_state_state;
  assign T30 = T25 & hit;
  assign hit = way_en != 4'h0;
  assign T31 = T32 ? io_way_en : way_en;
  assign T32 = state == 4'h4;
  assign T33 = T32 & T34;
  assign T34 = io_mshr_rdy ^ 1'h1;
  assign T35 = state == 4'h3;
  assign T36 = T37 & io_meta_read_ready;
  assign T37 = state == 4'h2;
  assign T38 = state == 4'h0;
  assign T39 = req_p_type == 2'h1;
  assign T40 = req_p_type == 2'h0;
  assign T41 = T46 ? 3'h1 : T42;
  assign T42 = T45 ? 3'h2 : T43;
  assign T43 = T44 ? 3'h3 : 3'h1;
  assign T44 = req_p_type == 2'h2;
  assign T45 = req_p_type == 2'h1;
  assign T46 = req_p_type == 2'h0;
  assign T47 = T48 == 2'h2;
  assign T48 = hit ? line_state_state : T49;
  assign T49 = 2'h0;
  assign io_wb_req_bits_client_xact_id = req_client_xact_id;
  assign T50 = T6 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_wb_req_bits_way_en = way_en;
  assign io_wb_req_bits_idx = T92;
  assign T92 = req_addr[3'h6:1'h0];
  assign T51 = T6 ? io_req_bits_addr : req_addr;
  assign io_wb_req_bits_tag = T52;
  assign T52 = req_addr >> 3'h7;
  assign io_wb_req_valid = T53;
  assign T53 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T54;
  assign T54 = T55;
  assign T55 = T60 ? 2'h0 : T56;
  assign T56 = T59 ? 2'h1 : T57;
  assign T57 = T58 ? line_state_state : line_state_state;
  assign T58 = req_p_type == 2'h2;
  assign T59 = req_p_type == 2'h1;
  assign T60 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T61;
  assign T61 = req_addr >> 3'h7;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T93;
  assign T93 = req_addr[3'h6:1'h0];
  assign io_meta_write_valid = T62;
  assign T62 = state == 4'h8;
  assign io_meta_read_bits_tag = T63;
  assign T63 = req_addr >> 3'h7;
  assign io_meta_read_bits_idx = T94;
  assign T94 = req_addr[3'h6:1'h0];
  assign io_meta_read_valid = T64;
  assign T64 = state == 4'h2;
  assign io_rep_bits_r_type = T65;
  assign T65 = T66;
  assign T66 = T79 ? T73 : T67;
  assign T67 = T72 ? 3'h4 : T68;
  assign T68 = T71 ? 3'h5 : T69;
  assign T69 = T70 ? 3'h6 : 3'h4;
  assign T70 = req_p_type == 2'h2;
  assign T71 = req_p_type == 2'h1;
  assign T72 = req_p_type == 2'h0;
  assign T73 = T78 ? 3'h1 : T74;
  assign T74 = T77 ? 3'h2 : T75;
  assign T75 = T76 ? 3'h3 : 3'h1;
  assign T76 = req_p_type == 2'h2;
  assign T77 = req_p_type == 2'h1;
  assign T78 = req_p_type == 2'h0;
  assign T79 = T80 == 2'h2;
  assign T80 = hit ? line_state_state : T81;
  assign T81 = 2'h0;
  assign io_rep_bits_data = T82;
  assign T82 = 136'h0;
  assign io_rep_bits_client_xact_id = T83;
  assign T83 = req_client_xact_id;
  assign io_rep_bits_addr = T84;
  assign T84 = req_addr;
  assign io_rep_valid = T85;
  assign T85 = T89 & T86;
  assign T86 = T87 ^ 1'h1;
  assign T87 = hit & T88;
  assign T88 = line_state_state == 2'h2;
  assign T89 = state == 4'h5;
  assign io_req_ready = T90;
  assign T90 = state == 4'h1;

  always @(posedge clk) begin
    if(T6) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(reset) begin
      state <= 4'h1;
    end else if(T38) begin
      state <= 4'h1;
    end else if(T6) begin
      state <= 4'h2;
    end else if(T36) begin
      state <= 4'h3;
    end else if(T35) begin
      state <= 4'h4;
    end else if(T33) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T30) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T23) begin
      state <= 4'h7;
    end else if(T21) begin
      state <= 4'h8;
    end else if(T19) begin
      state <= 4'h1;
    end
    if(T32) begin
      line_state_state <= io_line_state_state;
    end
    if(T32) begin
      way_en <= io_way_en;
    end
    if(T6) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T6) begin
      req_addr <= io_req_bits_addr;
    end
  end
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    input [18:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input [18:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[18:0] io_out_bits_tag,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[18:0] T0;
  wire T1;
  wire[6:0] T2;
  wire T3;
  wire T4;
  wire T5;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T0;
  assign T0 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T1 = chosen;
  assign io_out_bits_idx = T2;
  assign T2 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T3;
  assign T3 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T4;
  assign T4 = T5 & io_out_ready;
  assign T5 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [18:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [18:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[18:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[1:0] T0;
  wire T1;
  wire[18:0] T2;
  wire[3:0] T3;
  wire[6:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T0;
  assign T0 = T1 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T1 = chosen;
  assign io_out_bits_data_tag = T2;
  assign T2 = T1 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T3;
  assign T3 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T4;
  assign T4 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module LockingArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [135:0] io_in_1_bits_data,
    input  io_in_1_bits_uncached,
    input [1:0] io_in_1_bits_a_type,
    input [128:0] io_in_1_bits_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [135:0] io_in_0_bits_data,
    input  io_in_0_bits_uncached,
    input [1:0] io_in_0_bits_a_type,
    input [128:0] io_in_0_bits_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[135:0] io_out_bits_data,
    output io_out_bits_uncached,
    output[1:0] io_out_bits_a_type,
    output[128:0] io_out_bits_subblock,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T34;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  reg  locked;
  wire T35;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  reg [1:0] R17;
  wire[1:0] T36;
  wire[1:0] T18;
  wire[128:0] T19;
  wire T20;
  wire[1:0] T21;
  wire T22;
  wire[135:0] T23;
  wire[1:0] T24;
  wire[25:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R17 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T34 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T11 & T7;
  assign T7 = io_out_bits_uncached ? T8 : 1'h0;
  assign T8 = T10 | T9;
  assign T9 = 2'h2 == io_out_bits_a_type;
  assign T10 = 2'h1 == io_out_bits_a_type;
  assign T11 = io_out_ready & io_out_valid;
  assign T35 = reset ? 1'h0 : T12;
  assign T12 = T14 ? 1'h0 : T13;
  assign T13 = T4 ? 1'h1 : locked;
  assign T14 = T11 & T15;
  assign T15 = T16 == 2'h0;
  assign T16 = R17 + 2'h1;
  assign T36 = reset ? 2'h0 : T18;
  assign T18 = T6 ? T16 : R17;
  assign io_out_bits_subblock = T19;
  assign T19 = T20 ? io_in_1_bits_subblock : io_in_0_bits_subblock;
  assign T20 = chosen;
  assign io_out_bits_a_type = T21;
  assign T21 = T20 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_uncached = T22;
  assign T22 = T20 ? io_in_1_bits_uncached : io_in_0_bits_uncached;
  assign io_out_bits_data = T23;
  assign T23 = T20 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T24;
  assign T24 = T20 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T25;
  assign T25 = T20 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T26;
  assign T26 = T20 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = locked ? T29 : 1'h1;
  assign T29 = lockIdx == 1'h0;
  assign io_in_1_ready = T30;
  assign T30 = T31 & io_out_ready;
  assign T31 = locked ? T33 : T32;
  assign T32 = io_in_0_valid ^ 1'h1;
  assign T33 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T14) begin
      locked <= 1'h0;
    end else if(T4) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R17 <= 2'h0;
    end else if(T6) begin
      R17 <= T16;
    end
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[3:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_payload_manager_xact_id = T0;
  assign T0 = T1 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T1 = chosen;
  assign io_out_bits_header_dst = T2;
  assign T2 = T1 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T3;
  assign T3 = T1 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T4;
  assign T4 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [18:0] io_in_1_bits_tag,
    input [6:0] io_in_1_bits_idx,
    input [3:0] io_in_1_bits_way_en,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [18:0] io_in_0_bits_tag,
    input [6:0] io_in_0_bits_idx,
    input [3:0] io_in_0_bits_way_en,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[18:0] io_out_bits_tag,
    output[6:0] io_out_bits_idx,
    output[3:0] io_out_bits_way_en,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[2:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[3:0] T3;
  wire[6:0] T4;
  wire[18:0] T5;
  wire T6;
  wire T7;
  wire T8;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T0;
  assign T0 = T1 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T1 = chosen;
  assign io_out_bits_client_xact_id = T2;
  assign T2 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_way_en = T3;
  assign T3 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T4;
  assign T4 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_bits_tag = T5;
  assign T5 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_valid = T6;
  assign T6 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [3:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [7:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [3:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[3:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[7:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[4:0] T0;
  wire T1;
  wire[4:0] T2;
  wire[7:0] T3;
  wire[43:0] T4;
  wire T5;
  wire[3:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T0;
  assign T0 = T1 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T1 = chosen;
  assign io_out_bits_cmd = T2;
  assign T2 = T1 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T3;
  assign T3 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T4;
  assign T4 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T5;
  assign T5 = T1 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T6;
  assign T6 = T1 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T7;
  assign T7 = T1 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits = T0;
  assign T0 = T1 ? io_in_1_bits : io_in_0_bits;
  assign T1 = chosen;
  assign io_out_valid = T2;
  assign T2 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T3;
  assign T3 = T4 & io_out_ready;
  assign T4 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [3:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[3:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T29;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T30;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T31;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[67:0] T11;
  reg [67:0] ram [15:0];
  wire[67:0] T12;
  wire[67:0] T13;
  wire[67:0] T14;
  wire[61:0] T15;
  wire[9:0] T16;
  wire[51:0] T17;
  wire[5:0] T18;
  wire[4:0] T19;
  wire[4:0] T20;
  wire[7:0] T21;
  wire[43:0] T22;
  wire T23;
  wire[3:0] T24;
  wire T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T29 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T30 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T31 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_cmd, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_addr, io_enq_bits_tag};
  assign T18 = {io_enq_bits_kill, T19};
  assign T19 = {io_enq_bits_typ, io_enq_bits_phys};
  assign io_deq_bits_cmd = T20;
  assign T20 = T11[4'h9:3'h5];
  assign io_deq_bits_tag = T21;
  assign T21 = T11[5'h11:4'ha];
  assign io_deq_bits_addr = T22;
  assign T22 = T11[6'h3d:5'h12];
  assign io_deq_bits_phys = T23;
  assign T23 = T11[6'h3e:6'h3e];
  assign io_deq_bits_typ = T24;
  assign T24 = T11[7'h42:6'h3f];
  assign io_deq_bits_kill = T25;
  assign T25 = T11[7'h43:7'h43];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [3:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_idx_match,
    output[18:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[135:0] io_mem_req_bits_data,
    output io_mem_req_bits_uncached,
    output[1:0] io_mem_req_bits_a_type,
    output[128:0] io_mem_req_bits_subblock,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[135:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[3:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T0;
  wire can_finish;
  wire T1;
  reg [3:0] state;
  wire[3:0] T209;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire refill_done;
  wire T20;
  reg [1:0] refill_cnt;
  wire[1:0] T210;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire reply;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[3:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire wb_done;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire sec_rdy;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire idx_match;
  wire[6:0] T116;
  wire[6:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  reg [1:0] meta_hazard;
  wire[1:0] T211;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg [3:0] req_way_en;
  wire[3:0] T133;
  reg [18:0] req_old_meta_tag;
  wire[18:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[4:0] T138;
  wire[43:0] T212;
  wire[31:0] T139;
  wire[31:0] T140;
  wire[12:0] T141;
  wire[5:0] T142;
  wire T143;
  wire T144;
  wire[1:0] T145;
  reg [1:0] line_state_state;
  wire[1:0] T146;
  wire[1:0] T147;
  wire[1:0] T148;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T149;
  wire[1:0] T150;
  wire T151;
  wire T152;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire[1:0] meta_on_flush_state;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire[12:0] T166;
  wire[8:0] T167;
  wire[128:0] T168;
  wire[1:0] T169;
  reg [1:0] acquire_type;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[1:0] T213;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[135:0] T197;
  wire[1:0] T198;
  wire[25:0] T199;
  wire[25:0] T200;
  wire[25:0] T201;
  wire T202;
  wire T203;
  wire[18:0] T214;
  wire[30:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[3:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[3:0] ackq_io_deq_bits_payload_manager_xact_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    acquire_type = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_mem_finish_ready & can_finish;
  assign can_finish = T62 | T1;
  assign T1 = state == 4'h5;
  assign T209 = reset ? 4'h0 : T2;
  assign T2 = T60 ? T58 : T3;
  assign T3 = T56 ? 4'h4 : T4;
  assign T4 = T38 ? 4'h6 : T5;
  assign T5 = T37 ? 4'h2 : T6;
  assign T6 = T35 ? 4'h3 : T7;
  assign T7 = T33 ? 4'h4 : T8;
  assign T8 = T32 ? 4'h5 : T9;
  assign T9 = T19 ? 4'h6 : T10;
  assign T10 = T17 ? 4'h7 : T11;
  assign T11 = T16 ? 4'h8 : T12;
  assign T12 = T13 ? 4'h0 : state;
  assign T13 = T15 & T14;
  assign T14 = rpq_io_deq_valid ^ 1'h1;
  assign T15 = state == 4'h8;
  assign T16 = state == 4'h7;
  assign T17 = T18 & io_meta_write_ready;
  assign T18 = state == 4'h6;
  assign T19 = T31 & refill_done;
  assign refill_done = T25 & T20;
  assign T20 = refill_cnt == 2'h3;
  assign T210 = reset ? 2'h0 : T21;
  assign T21 = T24 ? 2'h0 : T22;
  assign T22 = T25 ? T23 : refill_cnt;
  assign T23 = refill_cnt + 2'h1;
  assign T24 = io_req_pri_val & io_req_pri_rdy;
  assign T25 = reply & T26;
  assign T26 = io_mem_grant_bits_payload_uncached ? 1'h0 : T27;
  assign T27 = T29 | T28;
  assign T28 = io_mem_grant_bits_payload_g_type == 2'h2;
  assign T29 = io_mem_grant_bits_payload_g_type == 2'h1;
  assign reply = io_mem_grant_valid & T30;
  assign T30 = io_mem_grant_bits_payload_client_xact_id == 2'h0;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & reply;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T55 & T39;
  assign T39 = T44 ? T43 : T40;
  assign T40 = T42 | T41;
  assign T41 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T42 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T43 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_cmd == 5'h6;
  assign T46 = T48 | T47;
  assign T47 = io_req_bits_cmd == 5'h3;
  assign T48 = T52 | T49;
  assign T49 = T51 | T50;
  assign T50 = io_req_bits_cmd == 5'h4;
  assign T51 = io_req_bits_cmd[2'h3:2'h3];
  assign T52 = T54 | T53;
  assign T53 = io_req_bits_cmd == 5'h7;
  assign T54 = io_req_bits_cmd == 5'h1;
  assign T55 = T24 & io_req_bits_tag_match;
  assign T56 = T55 & T57;
  assign T57 = T39 ^ 1'h1;
  assign T58 = T59 ? 4'h1 : 4'h3;
  assign T59 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T60 = T24 & T61;
  assign T61 = io_req_bits_tag_match ^ 1'h1;
  assign T62 = T64 | T63;
  assign T63 = state == 4'h4;
  assign T64 = state == 4'h0;
  assign T65 = T68 & T66;
  assign T66 = io_mem_grant_bits_payload_uncached | T67;
  assign T67 = io_mem_grant_bits_payload_g_type != 2'h0;
  assign T68 = wb_done | refill_done;
  assign wb_done = reply & T69;
  assign T69 = state == 4'h2;
  assign T70 = T75 ? 1'h0 : T71;
  assign T71 = T73 | T72;
  assign T72 = state == 4'h0;
  assign T73 = io_replay_ready & T74;
  assign T74 = state == 4'h8;
  assign T75 = io_meta_read_ready ^ 1'h1;
  assign T76 = T81 & T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = io_req_bits_cmd == 5'h3;
  assign T80 = io_req_bits_cmd == 5'h2;
  assign T81 = T118 | T82;
  assign T82 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T83;
  assign T83 = T111 | T84;
  assign T84 = T108 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T100 | T87;
  assign T87 = T89 & T88;
  assign T88 = io_mem_req_bits_a_type != 2'h1;
  assign T89 = T91 | T90;
  assign T90 = io_req_bits_cmd == 5'h6;
  assign T91 = T93 | T92;
  assign T92 = io_req_bits_cmd == 5'h3;
  assign T93 = T97 | T94;
  assign T94 = T96 | T95;
  assign T95 = io_req_bits_cmd == 5'h4;
  assign T96 = io_req_bits_cmd[2'h3:2'h3];
  assign T97 = T99 | T98;
  assign T98 = io_req_bits_cmd == 5'h7;
  assign T99 = io_req_bits_cmd == 5'h1;
  assign T100 = T101 & io_mem_req_bits_uncached;
  assign T101 = T105 | T102;
  assign T102 = T104 | T103;
  assign T103 = io_req_bits_cmd == 5'h4;
  assign T104 = io_req_bits_cmd[2'h3:2'h3];
  assign T105 = T107 | T106;
  assign T106 = io_req_bits_cmd == 5'h6;
  assign T107 = io_req_bits_cmd == 5'h0;
  assign T108 = T110 | T109;
  assign T109 = state == 4'h5;
  assign T110 = state == 4'h4;
  assign T111 = T113 | T112;
  assign T112 = state == 4'h3;
  assign T113 = T115 | T114;
  assign T114 = state == 4'h2;
  assign T115 = state == 4'h1;
  assign idx_match = req_idx == T116;
  assign T116 = io_req_bits_addr[4'hc:3'h6];
  assign req_idx = req_addr[4'hc:3'h6];
  assign T117 = T24 ? io_req_bits_addr : req_addr;
  assign T118 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T119;
  assign T119 = T132 | T120;
  assign T120 = T127 & T121;
  assign T121 = meta_hazard == 2'h0;
  assign T211 = reset ? 2'h0 : T122;
  assign T122 = T126 ? 2'h1 : T123;
  assign T123 = T125 ? T124 : meta_hazard;
  assign T124 = meta_hazard + 2'h1;
  assign T125 = meta_hazard != 2'h0;
  assign T126 = io_meta_write_ready & io_meta_write_valid;
  assign T127 = T129 & T128;
  assign T128 = state != 4'h3;
  assign T129 = T131 & T130;
  assign T130 = state != 4'h2;
  assign T131 = state != 4'h1;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h0;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T24 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T134 = T24 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T135;
  assign T135 = T136 & ackq_io_enq_ready;
  assign T136 = state == 4'h1;
  assign io_mem_finish_bits_payload_manager_xact_id = ackq_io_deq_bits_payload_manager_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T137;
  assign T137 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T138;
  assign T138 = T75 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T212;
  assign T212 = {12'h0, T139};
  assign T139 = T140;
  assign T140 = {io_tag, T141};
  assign T141 = {req_idx, T142};
  assign T142 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T143;
  assign T143 = T144 & rpq_io_deq_valid;
  assign T144 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T145;
  assign T145 = T161 ? meta_on_flush_state : line_state_state;
  assign T146 = T38 ? meta_on_hit_state : T147;
  assign T147 = T24 ? meta_on_flush_state : T148;
  assign T148 = T152 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T149;
  assign T149 = io_mem_grant_bits_payload_uncached ? 2'h0 : T150;
  assign T150 = T151 ? 2'h1 : 2'h2;
  assign T151 = io_mem_grant_bits_payload_g_type == 2'h1;
  assign T152 = T31 & reply;
  assign meta_on_hit_state = T153;
  assign T153 = T154 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign T154 = T158 | T155;
  assign T155 = T157 | T156;
  assign T156 = io_req_bits_cmd == 5'h4;
  assign T157 = io_req_bits_cmd[2'h3:2'h3];
  assign T158 = T160 | T159;
  assign T159 = io_req_bits_cmd == 5'h7;
  assign T160 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T161 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T162;
  assign T162 = T164 | T163;
  assign T163 = state == 4'h3;
  assign T164 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T165;
  assign T165 = state == 4'h8;
  assign io_mem_resp_data = {5{$random}};
  assign io_mem_resp_wmask = {1{$random}};
  assign io_mem_resp_addr = T166;
  assign T166 = T167 << 3'h4;
  assign T167 = {req_idx, refill_cnt};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_subblock = T168;
  assign T168 = 129'h0;
  assign io_mem_req_bits_a_type = T169;
  assign T169 = acquire_type;
  assign T170 = T24 ? T213 : T171;
  assign T171 = T184 ? T172 : acquire_type;
  assign T172 = T173 ? 2'h1 : io_mem_req_bits_a_type;
  assign T173 = T175 | T174;
  assign T174 = io_req_bits_cmd == 5'h6;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h3;
  assign T177 = T181 | T178;
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h4;
  assign T180 = io_req_bits_cmd[2'h3:2'h3];
  assign T181 = T183 | T182;
  assign T182 = io_req_bits_cmd == 5'h7;
  assign T183 = io_req_bits_cmd == 5'h1;
  assign T184 = io_req_sec_val & io_req_sec_rdy;
  assign T213 = {1'h0, T185};
  assign T185 = T187 | T186;
  assign T186 = io_req_bits_cmd == 5'h6;
  assign T187 = T189 | T188;
  assign T188 = io_req_bits_cmd == 5'h3;
  assign T189 = T193 | T190;
  assign T190 = T192 | T191;
  assign T191 = io_req_bits_cmd == 5'h4;
  assign T192 = io_req_bits_cmd[2'h3:2'h3];
  assign T193 = T195 | T194;
  assign T194 = io_req_bits_cmd == 5'h7;
  assign T195 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_uncached = T196;
  assign T196 = 1'h0;
  assign io_mem_req_bits_data = T197;
  assign T197 = 136'h0;
  assign io_mem_req_bits_client_xact_id = T198;
  assign T198 = 2'h0;
  assign io_mem_req_bits_addr = T199;
  assign T199 = T200;
  assign T200 = T201;
  assign T201 = {io_tag, req_idx};
  assign io_mem_req_valid = T202;
  assign T202 = T203 & ackq_io_enq_ready;
  assign T203 = state == 4'h4;
  assign io_tag = T214;
  assign T214 = T204[5'h12:1'h0];
  assign T204 = req_addr >> 4'hd;
  assign io_idx_match = T205;
  assign T205 = T206 & idx_match;
  assign T206 = state != 4'h0;
  assign io_req_sec_rdy = T207;
  assign T207 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T208;
  assign T208 = state == 4'h0;
  Queue_12 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T76 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T70 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_8 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T65 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( ackq_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ackq.io_enq_bits_header_src = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T60) begin
      state <= T58;
    end else if(T56) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T19) begin
      state <= 4'h6;
    end else if(T17) begin
      state <= 4'h7;
    end else if(T16) begin
      state <= 4'h8;
    end else if(T13) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T24) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T23;
    end
    if(T24) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T126) begin
      meta_hazard <= 2'h1;
    end else if(T125) begin
      meta_hazard <= T124;
    end
    if(T24) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T24) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T38) begin
      line_state_state <= meta_on_hit_state;
    end else if(T24) begin
      line_state_state <= meta_on_flush_state;
    end else if(T152) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T24) begin
      acquire_type <= T213;
    end else if(T184) begin
      acquire_type <= T172;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [3:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_idx_match,
    output[18:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[135:0] io_mem_req_bits_data,
    output io_mem_req_bits_uncached,
    output[1:0] io_mem_req_bits_a_type,
    output[128:0] io_mem_req_bits_subblock,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[135:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[3:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T0;
  wire can_finish;
  wire T1;
  reg [3:0] state;
  wire[3:0] T209;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire refill_done;
  wire T20;
  reg [1:0] refill_cnt;
  wire[1:0] T210;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire reply;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[3:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire wb_done;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire sec_rdy;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire idx_match;
  wire[6:0] T116;
  wire[6:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  reg [1:0] meta_hazard;
  wire[1:0] T211;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg [3:0] req_way_en;
  wire[3:0] T133;
  reg [18:0] req_old_meta_tag;
  wire[18:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[4:0] T138;
  wire[43:0] T212;
  wire[31:0] T139;
  wire[31:0] T140;
  wire[12:0] T141;
  wire[5:0] T142;
  wire T143;
  wire T144;
  wire[1:0] T145;
  reg [1:0] line_state_state;
  wire[1:0] T146;
  wire[1:0] T147;
  wire[1:0] T148;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T149;
  wire[1:0] T150;
  wire T151;
  wire T152;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire[1:0] meta_on_flush_state;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire[12:0] T166;
  wire[8:0] T167;
  wire[128:0] T168;
  wire[1:0] T169;
  reg [1:0] acquire_type;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[1:0] T213;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[135:0] T197;
  wire[1:0] T198;
  wire[25:0] T199;
  wire[25:0] T200;
  wire[25:0] T201;
  wire T202;
  wire T203;
  wire[18:0] T214;
  wire[30:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[3:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[3:0] ackq_io_deq_bits_payload_manager_xact_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    acquire_type = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_mem_finish_ready & can_finish;
  assign can_finish = T62 | T1;
  assign T1 = state == 4'h5;
  assign T209 = reset ? 4'h0 : T2;
  assign T2 = T60 ? T58 : T3;
  assign T3 = T56 ? 4'h4 : T4;
  assign T4 = T38 ? 4'h6 : T5;
  assign T5 = T37 ? 4'h2 : T6;
  assign T6 = T35 ? 4'h3 : T7;
  assign T7 = T33 ? 4'h4 : T8;
  assign T8 = T32 ? 4'h5 : T9;
  assign T9 = T19 ? 4'h6 : T10;
  assign T10 = T17 ? 4'h7 : T11;
  assign T11 = T16 ? 4'h8 : T12;
  assign T12 = T13 ? 4'h0 : state;
  assign T13 = T15 & T14;
  assign T14 = rpq_io_deq_valid ^ 1'h1;
  assign T15 = state == 4'h8;
  assign T16 = state == 4'h7;
  assign T17 = T18 & io_meta_write_ready;
  assign T18 = state == 4'h6;
  assign T19 = T31 & refill_done;
  assign refill_done = T25 & T20;
  assign T20 = refill_cnt == 2'h3;
  assign T210 = reset ? 2'h0 : T21;
  assign T21 = T24 ? 2'h0 : T22;
  assign T22 = T25 ? T23 : refill_cnt;
  assign T23 = refill_cnt + 2'h1;
  assign T24 = io_req_pri_val & io_req_pri_rdy;
  assign T25 = reply & T26;
  assign T26 = io_mem_grant_bits_payload_uncached ? 1'h0 : T27;
  assign T27 = T29 | T28;
  assign T28 = io_mem_grant_bits_payload_g_type == 2'h2;
  assign T29 = io_mem_grant_bits_payload_g_type == 2'h1;
  assign reply = io_mem_grant_valid & T30;
  assign T30 = io_mem_grant_bits_payload_client_xact_id == 2'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & reply;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T55 & T39;
  assign T39 = T44 ? T43 : T40;
  assign T40 = T42 | T41;
  assign T41 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T42 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T43 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_cmd == 5'h6;
  assign T46 = T48 | T47;
  assign T47 = io_req_bits_cmd == 5'h3;
  assign T48 = T52 | T49;
  assign T49 = T51 | T50;
  assign T50 = io_req_bits_cmd == 5'h4;
  assign T51 = io_req_bits_cmd[2'h3:2'h3];
  assign T52 = T54 | T53;
  assign T53 = io_req_bits_cmd == 5'h7;
  assign T54 = io_req_bits_cmd == 5'h1;
  assign T55 = T24 & io_req_bits_tag_match;
  assign T56 = T55 & T57;
  assign T57 = T39 ^ 1'h1;
  assign T58 = T59 ? 4'h1 : 4'h3;
  assign T59 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T60 = T24 & T61;
  assign T61 = io_req_bits_tag_match ^ 1'h1;
  assign T62 = T64 | T63;
  assign T63 = state == 4'h4;
  assign T64 = state == 4'h0;
  assign T65 = T68 & T66;
  assign T66 = io_mem_grant_bits_payload_uncached | T67;
  assign T67 = io_mem_grant_bits_payload_g_type != 2'h0;
  assign T68 = wb_done | refill_done;
  assign wb_done = reply & T69;
  assign T69 = state == 4'h2;
  assign T70 = T75 ? 1'h0 : T71;
  assign T71 = T73 | T72;
  assign T72 = state == 4'h0;
  assign T73 = io_replay_ready & T74;
  assign T74 = state == 4'h8;
  assign T75 = io_meta_read_ready ^ 1'h1;
  assign T76 = T81 & T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = io_req_bits_cmd == 5'h3;
  assign T80 = io_req_bits_cmd == 5'h2;
  assign T81 = T118 | T82;
  assign T82 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T83;
  assign T83 = T111 | T84;
  assign T84 = T108 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T100 | T87;
  assign T87 = T89 & T88;
  assign T88 = io_mem_req_bits_a_type != 2'h1;
  assign T89 = T91 | T90;
  assign T90 = io_req_bits_cmd == 5'h6;
  assign T91 = T93 | T92;
  assign T92 = io_req_bits_cmd == 5'h3;
  assign T93 = T97 | T94;
  assign T94 = T96 | T95;
  assign T95 = io_req_bits_cmd == 5'h4;
  assign T96 = io_req_bits_cmd[2'h3:2'h3];
  assign T97 = T99 | T98;
  assign T98 = io_req_bits_cmd == 5'h7;
  assign T99 = io_req_bits_cmd == 5'h1;
  assign T100 = T101 & io_mem_req_bits_uncached;
  assign T101 = T105 | T102;
  assign T102 = T104 | T103;
  assign T103 = io_req_bits_cmd == 5'h4;
  assign T104 = io_req_bits_cmd[2'h3:2'h3];
  assign T105 = T107 | T106;
  assign T106 = io_req_bits_cmd == 5'h6;
  assign T107 = io_req_bits_cmd == 5'h0;
  assign T108 = T110 | T109;
  assign T109 = state == 4'h5;
  assign T110 = state == 4'h4;
  assign T111 = T113 | T112;
  assign T112 = state == 4'h3;
  assign T113 = T115 | T114;
  assign T114 = state == 4'h2;
  assign T115 = state == 4'h1;
  assign idx_match = req_idx == T116;
  assign T116 = io_req_bits_addr[4'hc:3'h6];
  assign req_idx = req_addr[4'hc:3'h6];
  assign T117 = T24 ? io_req_bits_addr : req_addr;
  assign T118 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T119;
  assign T119 = T132 | T120;
  assign T120 = T127 & T121;
  assign T121 = meta_hazard == 2'h0;
  assign T211 = reset ? 2'h0 : T122;
  assign T122 = T126 ? 2'h1 : T123;
  assign T123 = T125 ? T124 : meta_hazard;
  assign T124 = meta_hazard + 2'h1;
  assign T125 = meta_hazard != 2'h0;
  assign T126 = io_meta_write_ready & io_meta_write_valid;
  assign T127 = T129 & T128;
  assign T128 = state != 4'h3;
  assign T129 = T131 & T130;
  assign T130 = state != 4'h2;
  assign T131 = state != 4'h1;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T24 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T134 = T24 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T135;
  assign T135 = T136 & ackq_io_enq_ready;
  assign T136 = state == 4'h1;
  assign io_mem_finish_bits_payload_manager_xact_id = ackq_io_deq_bits_payload_manager_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T137;
  assign T137 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T138;
  assign T138 = T75 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T212;
  assign T212 = {12'h0, T139};
  assign T139 = T140;
  assign T140 = {io_tag, T141};
  assign T141 = {req_idx, T142};
  assign T142 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T143;
  assign T143 = T144 & rpq_io_deq_valid;
  assign T144 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T145;
  assign T145 = T161 ? meta_on_flush_state : line_state_state;
  assign T146 = T38 ? meta_on_hit_state : T147;
  assign T147 = T24 ? meta_on_flush_state : T148;
  assign T148 = T152 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T149;
  assign T149 = io_mem_grant_bits_payload_uncached ? 2'h0 : T150;
  assign T150 = T151 ? 2'h1 : 2'h2;
  assign T151 = io_mem_grant_bits_payload_g_type == 2'h1;
  assign T152 = T31 & reply;
  assign meta_on_hit_state = T153;
  assign T153 = T154 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign T154 = T158 | T155;
  assign T155 = T157 | T156;
  assign T156 = io_req_bits_cmd == 5'h4;
  assign T157 = io_req_bits_cmd[2'h3:2'h3];
  assign T158 = T160 | T159;
  assign T159 = io_req_bits_cmd == 5'h7;
  assign T160 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T161 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T162;
  assign T162 = T164 | T163;
  assign T163 = state == 4'h3;
  assign T164 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T165;
  assign T165 = state == 4'h8;
  assign io_mem_resp_data = {5{$random}};
  assign io_mem_resp_wmask = {1{$random}};
  assign io_mem_resp_addr = T166;
  assign T166 = T167 << 3'h4;
  assign T167 = {req_idx, refill_cnt};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_subblock = T168;
  assign T168 = 129'h0;
  assign io_mem_req_bits_a_type = T169;
  assign T169 = acquire_type;
  assign T170 = T24 ? T213 : T171;
  assign T171 = T184 ? T172 : acquire_type;
  assign T172 = T173 ? 2'h1 : io_mem_req_bits_a_type;
  assign T173 = T175 | T174;
  assign T174 = io_req_bits_cmd == 5'h6;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h3;
  assign T177 = T181 | T178;
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h4;
  assign T180 = io_req_bits_cmd[2'h3:2'h3];
  assign T181 = T183 | T182;
  assign T182 = io_req_bits_cmd == 5'h7;
  assign T183 = io_req_bits_cmd == 5'h1;
  assign T184 = io_req_sec_val & io_req_sec_rdy;
  assign T213 = {1'h0, T185};
  assign T185 = T187 | T186;
  assign T186 = io_req_bits_cmd == 5'h6;
  assign T187 = T189 | T188;
  assign T188 = io_req_bits_cmd == 5'h3;
  assign T189 = T193 | T190;
  assign T190 = T192 | T191;
  assign T191 = io_req_bits_cmd == 5'h4;
  assign T192 = io_req_bits_cmd[2'h3:2'h3];
  assign T193 = T195 | T194;
  assign T194 = io_req_bits_cmd == 5'h7;
  assign T195 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_uncached = T196;
  assign T196 = 1'h0;
  assign io_mem_req_bits_data = T197;
  assign T197 = 136'h0;
  assign io_mem_req_bits_client_xact_id = T198;
  assign T198 = 2'h1;
  assign io_mem_req_bits_addr = T199;
  assign T199 = T200;
  assign T200 = T201;
  assign T201 = {io_tag, req_idx};
  assign io_mem_req_valid = T202;
  assign T202 = T203 & ackq_io_enq_ready;
  assign T203 = state == 4'h4;
  assign io_tag = T214;
  assign T214 = T204[5'h12:1'h0];
  assign T204 = req_addr >> 4'hd;
  assign io_idx_match = T205;
  assign T205 = T206 & idx_match;
  assign T206 = state != 4'h0;
  assign io_req_sec_rdy = T207;
  assign T207 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T208;
  assign T208 = state == 4'h0;
  Queue_12 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T76 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T70 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_8 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T65 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( ackq_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ackq.io_enq_bits_header_src = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T60) begin
      state <= T58;
    end else if(T56) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T19) begin
      state <= 4'h6;
    end else if(T17) begin
      state <= 4'h7;
    end else if(T16) begin
      state <= 4'h8;
    end else if(T13) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T24) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T23;
    end
    if(T24) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T126) begin
      meta_hazard <= 2'h1;
    end else if(T125) begin
      meta_hazard <= T124;
    end
    if(T24) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T24) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T38) begin
      line_state_state <= meta_on_hit_state;
    end else if(T24) begin
      line_state_state <= meta_on_flush_state;
    end else if(T152) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T24) begin
      acquire_type <= T213;
    end else if(T184) begin
      acquire_type <= T172;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input  io_req_bits_kill,
    input [3:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [63:0] io_req_bits_data,
    input  io_req_bits_tag_match,
    input [18:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input [3:0] io_req_bits_way_en,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[135:0] io_mem_req_bits_data,
    output io_mem_req_bits_uncached,
    output[1:0] io_mem_req_bits_a_type,
    output[128:0] io_mem_req_bits_subblock,
    output[3:0] io_mem_resp_way_en,
    output[12:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[135:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[6:0] io_meta_read_bits_idx,
    output[18:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[6:0] io_meta_write_bits_idx,
    output[3:0] io_meta_write_bits_way_en,
    output[18:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[3:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[63:0] io_replay_bits_data,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[18:0] io_wb_req_bits_tag,
    output[6:0] io_wb_req_bits_idx,
    output[3:0] io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire[4:0] T99;
  wire[4:0] T100;
  wire[4:0] T101;
  wire[4:0] T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire[4:0] T106;
  wire[4:0] T107;
  wire[4:0] T108;
  wire[4:0] T109;
  wire[4:0] T110;
  wire[4:0] T111;
  wire[4:0] T112;
  wire[4:0] T113;
  wire[4:0] T114;
  wire T115;
  wire[16:0] T0;
  wire[16:0] T1;
  reg [16:0] sdq_val;
  wire[16:0] T116;
  wire[31:0] T117;
  wire[31:0] T2;
  wire[31:0] T118;
  wire[31:0] T3;
  wire[31:0] T119;
  wire[16:0] T4;
  wire[16:0] T5;
  wire[16:0] T120;
  wire sdq_enq;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire[16:0] T14;
  wire[16:0] T15;
  wire[16:0] T16;
  wire[16:0] T17;
  wire[16:0] T18;
  wire[16:0] T19;
  wire[16:0] T20;
  wire[16:0] T21;
  wire[16:0] T22;
  wire[16:0] T23;
  wire[16:0] T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire[31:0] T51;
  wire[31:0] T52;
  wire[31:0] T121;
  wire[16:0] T53;
  wire[16:0] T122;
  wire free_sdq;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[31:0] T62;
  wire[31:0] T123;
  wire T63;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T64;
  wire tag_match;
  wire[30:0] T65;
  wire[30:0] T139;
  wire[18:0] T66;
  wire[18:0] T67;
  wire[18:0] tagList_1;
  wire idxMatch_1;
  wire[18:0] T68;
  wire[18:0] tagList_0;
  wire idxMatch_0;
  wire T69;
  wire sdq_rdy;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire idx_match;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire[63:0] T84;
  reg [63:0] sdq [16:0];
  wire[63:0] T85;
  wire T86;
  wire T87;
  wire[4:0] T88;
  reg [4:0] R89;
  wire[4:0] T90;
  wire[135:0] T91;
  wire[135:0] memRespMux_0_data;
  wire[135:0] memRespMux_1_data;
  wire T92;
  wire T140;
  wire[1:0] T93;
  wire[1:0] memRespMux_0_wmask;
  wire[1:0] memRespMux_1_wmask;
  wire[12:0] T94;
  wire[12:0] memRespMux_0_addr;
  wire[12:0] memRespMux_1_addr;
  wire[3:0] T95;
  wire[3:0] memRespMux_0_way_en;
  wire[3:0] memRespMux_1_way_en;
  wire T96;
  wire T97;
  wire pri_rdy;
  wire T98;
  wire sec_rdy;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[6:0] meta_read_arb_io_out_bits_idx;
  wire[18:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[6:0] meta_write_arb_io_out_bits_idx;
  wire[3:0] meta_write_arb_io_out_bits_way_en;
  wire[18:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr;
  wire[1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[135:0] mem_req_arb_io_out_bits_data;
  wire mem_req_arb_io_out_bits_uncached;
  wire[1:0] mem_req_arb_io_out_bits_a_type;
  wire[128:0] mem_req_arb_io_out_bits_subblock;
  wire mem_finish_arb_io_in_1_ready;
  wire mem_finish_arb_io_in_0_ready;
  wire mem_finish_arb_io_out_valid;
  wire[1:0] mem_finish_arb_io_out_bits_header_src;
  wire[1:0] mem_finish_arb_io_out_bits_header_dst;
  wire[3:0] mem_finish_arb_io_out_bits_payload_manager_xact_id;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[18:0] wb_req_arb_io_out_bits_tag;
  wire[6:0] wb_req_arb_io_out_bits_idx;
  wire[3:0] wb_req_arb_io_out_bits_way_en;
  wire[1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire replay_arb_io_out_bits_kill;
  wire[3:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_phys;
  wire[43:0] replay_arb_io_out_bits_addr;
  wire[7:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire MSHR_0_io_req_pri_rdy;
  wire MSHR_0_io_req_sec_rdy;
  wire MSHR_0_io_idx_match;
  wire[18:0] MSHR_0_io_tag;
  wire MSHR_0_io_mem_req_valid;
  wire[25:0] MSHR_0_io_mem_req_bits_addr;
  wire[1:0] MSHR_0_io_mem_req_bits_client_xact_id;
  wire[135:0] MSHR_0_io_mem_req_bits_data;
  wire MSHR_0_io_mem_req_bits_uncached;
  wire[1:0] MSHR_0_io_mem_req_bits_a_type;
  wire[128:0] MSHR_0_io_mem_req_bits_subblock;
  wire[3:0] MSHR_0_io_mem_resp_way_en;
  wire[12:0] MSHR_0_io_mem_resp_addr;
  wire[1:0] MSHR_0_io_mem_resp_wmask;
  wire[135:0] MSHR_0_io_mem_resp_data;
  wire MSHR_0_io_meta_read_valid;
  wire[6:0] MSHR_0_io_meta_read_bits_idx;
  wire[18:0] MSHR_0_io_meta_read_bits_tag;
  wire MSHR_0_io_meta_write_valid;
  wire[6:0] MSHR_0_io_meta_write_bits_idx;
  wire[3:0] MSHR_0_io_meta_write_bits_way_en;
  wire[18:0] MSHR_0_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_0_io_meta_write_bits_data_coh_state;
  wire MSHR_0_io_replay_valid;
  wire MSHR_0_io_replay_bits_kill;
  wire[3:0] MSHR_0_io_replay_bits_typ;
  wire MSHR_0_io_replay_bits_phys;
  wire[43:0] MSHR_0_io_replay_bits_addr;
  wire[7:0] MSHR_0_io_replay_bits_tag;
  wire[4:0] MSHR_0_io_replay_bits_cmd;
  wire[4:0] MSHR_0_io_replay_bits_sdq_id;
  wire MSHR_0_io_mem_finish_valid;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_dst;
  wire[3:0] MSHR_0_io_mem_finish_bits_payload_manager_xact_id;
  wire MSHR_0_io_wb_req_valid;
  wire[18:0] MSHR_0_io_wb_req_bits_tag;
  wire[6:0] MSHR_0_io_wb_req_bits_idx;
  wire[3:0] MSHR_0_io_wb_req_bits_way_en;
  wire[1:0] MSHR_0_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_0_io_wb_req_bits_r_type;
  wire MSHR_0_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[18:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr;
  wire[1:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[135:0] MSHR_1_io_mem_req_bits_data;
  wire MSHR_1_io_mem_req_bits_uncached;
  wire[1:0] MSHR_1_io_mem_req_bits_a_type;
  wire[128:0] MSHR_1_io_mem_req_bits_subblock;
  wire[3:0] MSHR_1_io_mem_resp_way_en;
  wire[12:0] MSHR_1_io_mem_resp_addr;
  wire[1:0] MSHR_1_io_mem_resp_wmask;
  wire[135:0] MSHR_1_io_mem_resp_data;
  wire MSHR_1_io_meta_read_valid;
  wire[6:0] MSHR_1_io_meta_read_bits_idx;
  wire[18:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[6:0] MSHR_1_io_meta_write_bits_idx;
  wire[3:0] MSHR_1_io_meta_write_bits_way_en;
  wire[18:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire MSHR_1_io_replay_bits_kill;
  wire[3:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_phys;
  wire[43:0] MSHR_1_io_replay_bits_addr;
  wire[7:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_mem_finish_valid;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_dst;
  wire[3:0] MSHR_1_io_mem_finish_bits_payload_manager_xact_id;
  wire MSHR_1_io_wb_req_valid;
  wire[18:0] MSHR_1_io_wb_req_bits_tag;
  wire[6:0] MSHR_1_io_wb_req_bits_idx;
  wire[3:0] MSHR_1_io_wb_req_bits_way_en;
  wire[1:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R89 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T99 = T138 ? 1'h0 : T100;
  assign T100 = T137 ? 1'h1 : T101;
  assign T101 = T136 ? 2'h2 : T102;
  assign T102 = T135 ? 2'h3 : T103;
  assign T103 = T134 ? 3'h4 : T104;
  assign T104 = T133 ? 3'h5 : T105;
  assign T105 = T132 ? 3'h6 : T106;
  assign T106 = T131 ? 3'h7 : T107;
  assign T107 = T130 ? 4'h8 : T108;
  assign T108 = T129 ? 4'h9 : T109;
  assign T109 = T128 ? 4'ha : T110;
  assign T110 = T127 ? 4'hb : T111;
  assign T111 = T126 ? 4'hc : T112;
  assign T112 = T125 ? 4'hd : T113;
  assign T113 = T124 ? 4'he : T114;
  assign T114 = T115 ? 4'hf : 5'h10;
  assign T115 = T0[4'hf:4'hf];
  assign T0 = ~ T1;
  assign T1 = sdq_val[5'h10:1'h0];
  assign T116 = T117[5'h10:1'h0];
  assign T117 = reset ? 32'h0 : T2;
  assign T2 = T63 ? T3 : T118;
  assign T118 = {15'h0, sdq_val};
  assign T3 = T50 | T119;
  assign T119 = {15'h0, T4};
  assign T4 = T14 & T5;
  assign T5 = 17'h0 - T120;
  assign T120 = {16'h0, sdq_enq};
  assign sdq_enq = T13 & T6;
  assign T6 = T10 | T7;
  assign T7 = T9 | T8;
  assign T8 = io_req_bits_cmd == 5'h4;
  assign T9 = io_req_bits_cmd[2'h3:2'h3];
  assign T10 = T12 | T11;
  assign T11 = io_req_bits_cmd == 5'h7;
  assign T12 = io_req_bits_cmd == 5'h1;
  assign T13 = io_req_valid & io_req_ready;
  assign T14 = T49 ? 17'h1 : T15;
  assign T15 = T48 ? 17'h2 : T16;
  assign T16 = T47 ? 17'h4 : T17;
  assign T17 = T46 ? 17'h8 : T18;
  assign T18 = T45 ? 17'h10 : T19;
  assign T19 = T44 ? 17'h20 : T20;
  assign T20 = T43 ? 17'h40 : T21;
  assign T21 = T42 ? 17'h80 : T22;
  assign T22 = T41 ? 17'h100 : T23;
  assign T23 = T40 ? 17'h200 : T24;
  assign T24 = T39 ? 17'h400 : T25;
  assign T25 = T38 ? 17'h800 : T26;
  assign T26 = T37 ? 17'h1000 : T27;
  assign T27 = T36 ? 17'h2000 : T28;
  assign T28 = T35 ? 17'h4000 : T29;
  assign T29 = T34 ? 17'h8000 : T30;
  assign T30 = T31 ? 17'h10000 : 17'h0;
  assign T31 = T32[5'h10:5'h10];
  assign T32 = ~ T33;
  assign T33 = sdq_val[5'h10:1'h0];
  assign T34 = T32[4'hf:4'hf];
  assign T35 = T32[4'he:4'he];
  assign T36 = T32[4'hd:4'hd];
  assign T37 = T32[4'hc:4'hc];
  assign T38 = T32[4'hb:4'hb];
  assign T39 = T32[4'ha:4'ha];
  assign T40 = T32[4'h9:4'h9];
  assign T41 = T32[4'h8:4'h8];
  assign T42 = T32[3'h7:3'h7];
  assign T43 = T32[3'h6:3'h6];
  assign T44 = T32[3'h5:3'h5];
  assign T45 = T32[3'h4:3'h4];
  assign T46 = T32[2'h3:2'h3];
  assign T47 = T32[2'h2:2'h2];
  assign T48 = T32[1'h1:1'h1];
  assign T49 = T32[1'h0:1'h0];
  assign T50 = T123 & T51;
  assign T51 = ~ T52;
  assign T52 = T62 & T121;
  assign T121 = {15'h0, T53};
  assign T53 = 17'h0 - T122;
  assign T122 = {16'h0, free_sdq};
  assign free_sdq = T61 & T54;
  assign T54 = T58 | T55;
  assign T55 = T57 | T56;
  assign T56 = io_replay_bits_cmd == 5'h4;
  assign T57 = io_replay_bits_cmd[2'h3:2'h3];
  assign T58 = T60 | T59;
  assign T59 = io_replay_bits_cmd == 5'h7;
  assign T60 = io_replay_bits_cmd == 5'h1;
  assign T61 = io_replay_ready & io_replay_valid;
  assign T62 = 1'h1 << replay_arb_io_out_bits_sdq_id;
  assign T123 = {15'h0, sdq_val};
  assign T63 = io_replay_valid | sdq_enq;
  assign T124 = T0[4'he:4'he];
  assign T125 = T0[4'hd:4'hd];
  assign T126 = T0[4'hc:4'hc];
  assign T127 = T0[4'hb:4'hb];
  assign T128 = T0[4'ha:4'ha];
  assign T129 = T0[4'h9:4'h9];
  assign T130 = T0[4'h8:4'h8];
  assign T131 = T0[3'h7:3'h7];
  assign T132 = T0[3'h6:3'h6];
  assign T133 = T0[3'h5:3'h5];
  assign T134 = T0[3'h4:3'h4];
  assign T135 = T0[2'h3:2'h3];
  assign T136 = T0[2'h2:2'h2];
  assign T137 = T0[1'h1:1'h1];
  assign T138 = T0[1'h0:1'h0];
  assign T64 = T69 & tag_match;
  assign tag_match = T139 == T65;
  assign T65 = io_req_bits_addr >> 4'hd;
  assign T139 = {12'h0, T66};
  assign T66 = T68 | T67;
  assign T67 = idxMatch_1 ? tagList_1 : 19'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T68 = idxMatch_0 ? tagList_0 : 19'h0;
  assign tagList_0 = MSHR_0_io_tag;
  assign idxMatch_0 = MSHR_0_io_idx_match;
  assign T69 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T70 ^ 1'h1;
  assign T70 = sdq_val == 17'h1ffff;
  assign T71 = T72 & tag_match;
  assign T72 = io_req_valid & sdq_rdy;
  assign T73 = T75 & T74;
  assign T74 = idx_match ^ 1'h1;
  assign idx_match = MSHR_0_io_idx_match | MSHR_1_io_idx_match;
  assign T75 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T76;
  assign T76 = T79 ? 1'h0 : T77;
  assign T77 = T78 == 1'h0;
  assign T78 = MSHR_0_io_req_pri_rdy ^ 1'h1;
  assign T79 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T80;
  assign T80 = T83 ? 1'h0 : T81;
  assign T81 = T82 == 1'h0;
  assign T82 = MSHR_0_io_probe_rdy ^ 1'h1;
  assign T83 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_idx = wb_req_arb_io_out_bits_idx;
  assign io_wb_req_bits_tag = wb_req_arb_io_out_bits_tag;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_mem_finish_bits_payload_manager_xact_id = mem_finish_arb_io_out_bits_payload_manager_xact_id;
  assign io_mem_finish_bits_header_dst = mem_finish_arb_io_out_bits_header_dst;
  assign io_mem_finish_bits_header_src = mem_finish_arb_io_out_bits_header_src;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_replay_bits_data = T84;
  assign T84 = sdq[R89];
  assign T86 = sdq_enq & T87;
  assign T87 = T88 < 5'h11;
  assign T88 = T99[3'h4:1'h0];
  assign T90 = free_sdq ? replay_arb_io_out_bits_sdq_id : R89;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_mem_resp_data = T91;
  assign T91 = T92 ? memRespMux_1_data : memRespMux_0_data;
  assign memRespMux_0_data = MSHR_0_io_mem_resp_data;
  assign memRespMux_1_data = MSHR_1_io_mem_resp_data;
  assign T92 = T140;
  assign T140 = io_mem_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_mem_resp_wmask = T93;
  assign T93 = T92 ? memRespMux_1_wmask : memRespMux_0_wmask;
  assign memRespMux_0_wmask = MSHR_0_io_mem_resp_wmask;
  assign memRespMux_1_wmask = MSHR_1_io_mem_resp_wmask;
  assign io_mem_resp_addr = T94;
  assign T94 = T92 ? memRespMux_1_addr : memRespMux_0_addr;
  assign memRespMux_0_addr = MSHR_0_io_mem_resp_addr;
  assign memRespMux_1_addr = MSHR_1_io_mem_resp_addr;
  assign io_mem_resp_way_en = T95;
  assign T95 = T92 ? memRespMux_1_way_en : memRespMux_0_way_en;
  assign memRespMux_0_way_en = MSHR_0_io_mem_resp_way_en;
  assign memRespMux_1_way_en = MSHR_1_io_mem_resp_way_en;
  assign io_mem_req_bits_subblock = mem_req_arb_io_out_bits_subblock;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_uncached = mem_req_arb_io_out_bits_uncached;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr = mem_req_arb_io_out_bits_addr;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T96;
  assign T96 = T97 & sdq_rdy;
  assign T97 = idx_match ? T98 : pri_rdy;
  assign pri_rdy = MSHR_0_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T98 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_0_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_5 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  LockingArbiter_1 mem_req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_in_1_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_in_1_bits_uncached( MSHR_1_io_mem_req_bits_uncached ),
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_in_1_bits_subblock( MSHR_1_io_mem_req_bits_subblock ),
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_req_valid ),
       .io_in_0_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       .io_in_0_bits_data( MSHR_0_io_mem_req_bits_data ),
       .io_in_0_bits_uncached( MSHR_0_io_mem_req_bits_uncached ),
       .io_in_0_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       .io_in_0_bits_subblock( MSHR_0_io_mem_req_bits_subblock ),
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr( mem_req_arb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_uncached( mem_req_arb_io_out_bits_uncached ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_subblock( mem_req_arb_io_out_bits_subblock )
       //.io_chosen(  )
  );
  Arbiter_6 mem_finish_arb(
       .io_in_1_ready( mem_finish_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_finish_valid ),
       .io_in_1_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_in_1_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( MSHR_1_io_mem_finish_bits_payload_manager_xact_id ),
       .io_in_0_ready( mem_finish_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_finish_valid ),
       .io_in_0_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_in_0_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( MSHR_0_io_mem_finish_bits_payload_manager_xact_id ),
       .io_out_ready( io_mem_finish_ready ),
       .io_out_valid( mem_finish_arb_io_out_valid ),
       .io_out_bits_header_src( mem_finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( mem_finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( mem_finish_arb_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_wb_req_valid ),
       .io_in_0_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_tag( wb_req_arb_io_out_bits_tag ),
       .io_out_bits_idx( wb_req_arb_io_out_bits_idx ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  Arbiter_7 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_replay_valid ),
       .io_in_0_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_in_0_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_in_0_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_in_0_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_in_0_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_in_0_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_8 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T73 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  MSHR_0 MSHR_0(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_0_io_req_pri_rdy ),
       .io_req_sec_val( T71 ),
       .io_req_sec_rdy( MSHR_0_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_sdq_id( T99 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_0_io_idx_match ),
       .io_tag( MSHR_0_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_0_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( MSHR_0_io_mem_req_bits_data ),
       .io_mem_req_bits_uncached( MSHR_0_io_mem_req_bits_uncached ),
       .io_mem_req_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       .io_mem_req_bits_subblock( MSHR_0_io_mem_req_bits_subblock ),
       .io_mem_resp_way_en( MSHR_0_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_0_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_0_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_0_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_0_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_0_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_0_io_replay_valid ),
       .io_replay_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_0_ready ),
       .io_mem_finish_valid( MSHR_0_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( MSHR_0_io_mem_finish_bits_payload_manager_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_0_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_0_io_probe_rdy )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MSHR_0.io_mem_resp_wmask = {1{$random}};
    assign MSHR_0.io_mem_resp_data = {5{$random}};
// synthesis translate_on
`endif
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T64 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_sdq_id( T99 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_mem_req_bits_uncached( MSHR_1_io_mem_req_bits_uncached ),
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_mem_req_bits_subblock( MSHR_1_io_mem_req_bits_subblock ),
       .io_mem_resp_way_en( MSHR_1_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_1_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_1_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_1_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_1_ready ),
       .io_mem_finish_valid( MSHR_1_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( MSHR_1_io_mem_finish_bits_payload_manager_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MSHR_1.io_mem_resp_wmask = {1{$random}};
    assign MSHR_1.io_mem_resp_data = {5{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    sdq_val <= T116;
    if (T86)
      sdq[T99] <= io_req_bits_data;
    if(free_sdq) begin
      R89 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [6:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [6:0] io_write_bits_idx,
    input [3:0] io_write_bits_way_en,
    input [18:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[18:0] io_resp_3_tag,
    output[1:0] io_resp_3_coh_state,
    output[18:0] io_resp_2_tag,
    output[1:0] io_resp_2_coh_state,
    output[18:0] io_resp_1_tag,
    output[1:0] io_resp_1_coh_state,
    output[18:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[20:0] T1;
  wire[83:0] tags;
  wire[83:0] T2;
  wire[83:0] T3;
  wire[83:0] T4;
  wire[41:0] T5;
  wire[20:0] T6;
  wire[20:0] T40;
  wire T7;
  wire[3:0] wmask;
  wire rst;
  reg [7:0] rst_cnt;
  wire[7:0] T41;
  wire[7:0] T8;
  wire[7:0] T9;
  wire[20:0] T10;
  wire[20:0] T42;
  wire T11;
  wire[41:0] T12;
  wire[20:0] T13;
  wire[20:0] T43;
  wire T14;
  wire[20:0] T15;
  wire[20:0] T44;
  wire T16;
  wire[83:0] T17;
  wire[41:0] T18;
  wire[20:0] wdata;
  wire[20:0] T19;
  wire[1:0] T20;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T21;
  wire[18:0] T22;
  wire[18:0] rstVal_tag;
  wire T23;
  wire[6:0] T45;
  wire[7:0] waddr;
  wire[7:0] T46;
  reg [6:0] R24;
  wire[6:0] T25;
  wire[18:0] T26;
  wire[1:0] T27;
  wire[20:0] T28;
  wire[18:0] T29;
  wire[1:0] T30;
  wire[20:0] T31;
  wire[18:0] T32;
  wire[1:0] T33;
  wire[20:0] T34;
  wire[18:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R24 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = tags[5'h14:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T45),
    .W0E(T23),
    .W0I(T17),
    .W0M(T3),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(tags)
  );
  assign T3 = T4;
  assign T4 = {T12, T5};
  assign T5 = {T10, T6};
  assign T6 = 21'h0 - T40;
  assign T40 = {20'h0, T7};
  assign T7 = wmask[1'h0:1'h0];
  assign wmask = rst ? 4'hf : io_write_bits_way_en;
  assign rst = rst_cnt < 8'h80;
  assign T41 = reset ? 8'h0 : T8;
  assign T8 = rst ? T9 : rst_cnt;
  assign T9 = rst_cnt + 8'h1;
  assign T10 = 21'h0 - T42;
  assign T42 = {20'h0, T11};
  assign T11 = wmask[1'h1:1'h1];
  assign T12 = {T15, T13};
  assign T13 = 21'h0 - T43;
  assign T43 = {20'h0, T14};
  assign T14 = wmask[2'h2:2'h2];
  assign T15 = 21'h0 - T44;
  assign T44 = {20'h0, T16};
  assign T16 = wmask[2'h3:2'h3];
  assign T17 = {T18, T18};
  assign T18 = {wdata, wdata};
  assign wdata = T19;
  assign T19 = {T22, T20};
  assign T20 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T21;
  assign T21 = 2'h0;
  assign T22 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 19'h0;
  assign T23 = rst | io_write_valid;
  assign T45 = waddr[3'h6:1'h0];
  assign waddr = rst ? rst_cnt : T46;
  assign T46 = {1'h0, io_write_bits_idx};
  assign T25 = io_read_valid ? io_read_bits_idx : R24;
  assign io_resp_0_tag = T26;
  assign T26 = T1[5'h14:2'h2];
  assign io_resp_1_coh_state = T27;
  assign T27 = T28[1'h1:1'h0];
  assign T28 = tags[6'h29:5'h15];
  assign io_resp_1_tag = T29;
  assign T29 = T28[5'h14:2'h2];
  assign io_resp_2_coh_state = T30;
  assign T30 = T31[1'h1:1'h0];
  assign T31 = tags[6'h3e:6'h2a];
  assign io_resp_2_tag = T32;
  assign T32 = T31[5'h14:2'h2];
  assign io_resp_3_coh_state = T33;
  assign T33 = T34[1'h1:1'h0];
  assign T34 = tags[7'h53:6'h3f];
  assign io_resp_3_tag = T35;
  assign T35 = T34[5'h14:2'h2];
  assign io_write_ready = T36;
  assign T36 = rst ^ 1'h1;
  assign io_read_ready = T37;
  assign T37 = T39 & T38;
  assign T38 = io_write_valid ^ 1'h1;
  assign T39 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 8'h0;
    end else if(rst) begin
      rst_cnt <= T9;
    end
    if(io_read_valid) begin
      R24 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [6:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [6:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [6:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [6:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [6:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[6:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire[6:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[6:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T3;
  assign T3 = T11 ? io_in_4_bits_idx : T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = chosen;
  assign T8 = T9 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign T11 = T7[2'h2:2'h2];
  assign io_out_valid = T12;
  assign T12 = T19 ? io_in_4_valid : T13;
  assign T13 = T18 ? T16 : T14;
  assign T14 = T15 ? io_in_1_valid : io_in_0_valid;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T17 ? io_in_3_valid : io_in_2_valid;
  assign T17 = T7[1'h0:1'h0];
  assign T18 = T7[1'h1:1'h1];
  assign T19 = T7[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = T28 | io_in_2_valid;
  assign T28 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T32 | io_in_3_valid;
  assign T32 = T33 | io_in_2_valid;
  assign T33 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input [3:0] io_read_bits_way_en,
    input [12:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input [3:0] io_write_bits_way_en,
    input [12:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [135:0] io_write_bits_data,
    output[135:0] io_resp_3,
    output[135:0] io_resp_2,
    output[135:0] io_resp_1,
    output[135:0] io_resp_0
);

  wire[135:0] T0;
  wire[135:0] T1;
  wire[67:0] T2;
  wire[67:0] T3;
  wire[135:0] T4;
  wire[135:0] T5;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire[8:0] raddr;
  wire[135:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[67:0] T10;
  wire[67:0] T116;
  wire T11;
  wire[1:0] T12;
  wire[67:0] T13;
  wire[67:0] T117;
  wire T14;
  wire[135:0] T15;
  wire[67:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[8:0] waddr;
  reg [8:0] R21;
  wire[8:0] T22;
  wire T26;
  wire T27;
  reg [12:0] R28;
  wire[12:0] T29;
  wire[67:0] T30;
  wire[135:0] T31;
  wire[135:0] T32;
  wire T49;
  wire T50;
  wire[135:0] T34;
  wire[135:0] T35;
  wire[135:0] T36;
  wire[67:0] T37;
  wire[67:0] T118;
  wire T38;
  wire[67:0] T39;
  wire[67:0] T119;
  wire T40;
  wire[135:0] T41;
  wire[67:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg [8:0] R47;
  wire[8:0] T48;
  wire[135:0] T51;
  wire[135:0] T52;
  wire[67:0] T53;
  wire[67:0] T54;
  wire T55;
  wire T56;
  wire[67:0] T57;
  wire[135:0] T58;
  wire[135:0] T59;
  wire[67:0] T60;
  wire[67:0] T61;
  wire[135:0] T62;
  wire[135:0] T63;
  wire T81;
  wire T82;
  wire[1:0] T83;
  wire[135:0] T65;
  wire[135:0] T66;
  wire[135:0] T67;
  wire[67:0] T68;
  wire[67:0] T120;
  wire T69;
  wire[1:0] T70;
  wire[67:0] T71;
  wire[67:0] T121;
  wire T72;
  wire[135:0] T73;
  wire[67:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [8:0] R79;
  wire[8:0] T80;
  wire T84;
  wire T85;
  reg [12:0] R86;
  wire[12:0] T87;
  wire[67:0] T88;
  wire[135:0] T89;
  wire[135:0] T90;
  wire T107;
  wire T108;
  wire[135:0] T92;
  wire[135:0] T93;
  wire[135:0] T94;
  wire[67:0] T95;
  wire[67:0] T122;
  wire T96;
  wire[67:0] T97;
  wire[67:0] T123;
  wire T98;
  wire[135:0] T99;
  wire[67:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg [8:0] R105;
  wire[8:0] T106;
  wire[135:0] T109;
  wire[135:0] T110;
  wire[67:0] T111;
  wire[67:0] T112;
  wire T113;
  wire T114;
  wire[67:0] T115;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R21 = {1{$random}};
    R28 = {1{$random}};
    R47 = {1{$random}};
    R79 = {1{$random}};
    R86 = {1{$random}};
    R105 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0 = T0;
  assign T0 = T1;
  assign T1 = {T30, T2};
  assign T2 = T26 ? T30 : T3;
  assign T3 = T4[7'h43:1'h0];
  assign T4 = T5;
  assign T23 = T24 & io_read_valid;
  assign T24 = T25 != 2'h0;
  assign T25 = io_read_bits_way_en[1'h1:1'h0];
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T6 T6 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T17),
    .W0I(T15),
    .W0M(T8),
    .R1A(raddr),
    .R1E(T23),
    .R1O(T5)
  );
  assign T8 = T9;
  assign T9 = {T13, T10};
  assign T10 = 68'h0 - T116;
  assign T116 = {67'h0, T11};
  assign T11 = T12[1'h0:1'h0];
  assign T12 = io_write_bits_way_en[1'h1:1'h0];
  assign T13 = 68'h0 - T117;
  assign T117 = {67'h0, T14};
  assign T14 = T12[1'h1:1'h1];
  assign T15 = {T16, T16};
  assign T16 = io_write_bits_data[7'h43:1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_write_bits_wmask[1'h0:1'h0];
  assign T19 = T20 & io_write_valid;
  assign T20 = T12 != 2'h0;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T22 = T23 ? raddr : R21;
  assign T26 = T27;
  assign T27 = R28[2'h3:2'h3];
  assign T29 = io_read_valid ? io_read_bits_addr : R28;
  assign T30 = T31[7'h43:1'h0];
  assign T31 = T32;
  assign T49 = T50 & io_read_valid;
  assign T50 = T25 != 2'h0;
  DataArray_T6 T33 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T43),
    .W0I(T41),
    .W0M(T35),
    .R1A(raddr),
    .R1E(T49),
    .R1O(T32)
  );
  assign T35 = T36;
  assign T36 = {T39, T37};
  assign T37 = 68'h0 - T118;
  assign T118 = {67'h0, T38};
  assign T38 = T12[1'h0:1'h0];
  assign T39 = 68'h0 - T119;
  assign T119 = {67'h0, T40};
  assign T40 = T12[1'h1:1'h1];
  assign T41 = {T42, T42};
  assign T42 = io_write_bits_data[8'h87:7'h44];
  assign T43 = T45 & T44;
  assign T44 = io_write_bits_wmask[1'h1:1'h1];
  assign T45 = T46 & io_write_valid;
  assign T46 = T12 != 2'h0;
  assign T48 = T49 ? raddr : R47;
  assign io_resp_1 = T51;
  assign T51 = T52;
  assign T52 = {T57, T53};
  assign T53 = T55 ? T57 : T54;
  assign T54 = T4[8'h87:7'h44];
  assign T55 = T56;
  assign T56 = R28[2'h3:2'h3];
  assign T57 = T31[8'h87:7'h44];
  assign io_resp_2 = T58;
  assign T58 = T59;
  assign T59 = {T88, T60};
  assign T60 = T84 ? T88 : T61;
  assign T61 = T62[7'h43:1'h0];
  assign T62 = T63;
  assign T81 = T82 & io_read_valid;
  assign T82 = T83 != 2'h0;
  assign T83 = io_read_bits_way_en[2'h3:2'h2];
  DataArray_T6 T64 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T75),
    .W0I(T73),
    .W0M(T66),
    .R1A(raddr),
    .R1E(T81),
    .R1O(T63)
  );
  assign T66 = T67;
  assign T67 = {T71, T68};
  assign T68 = 68'h0 - T120;
  assign T120 = {67'h0, T69};
  assign T69 = T70[1'h0:1'h0];
  assign T70 = io_write_bits_way_en[2'h3:2'h2];
  assign T71 = 68'h0 - T121;
  assign T121 = {67'h0, T72};
  assign T72 = T70[1'h1:1'h1];
  assign T73 = {T74, T74};
  assign T74 = io_write_bits_data[7'h43:1'h0];
  assign T75 = T77 & T76;
  assign T76 = io_write_bits_wmask[1'h0:1'h0];
  assign T77 = T78 & io_write_valid;
  assign T78 = T70 != 2'h0;
  assign T80 = T81 ? raddr : R79;
  assign T84 = T85;
  assign T85 = R86[2'h3:2'h3];
  assign T87 = io_read_valid ? io_read_bits_addr : R86;
  assign T88 = T89[7'h43:1'h0];
  assign T89 = T90;
  assign T107 = T108 & io_read_valid;
  assign T108 = T83 != 2'h0;
  DataArray_T6 T91 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T101),
    .W0I(T99),
    .W0M(T93),
    .R1A(raddr),
    .R1E(T107),
    .R1O(T90)
  );
  assign T93 = T94;
  assign T94 = {T97, T95};
  assign T95 = 68'h0 - T122;
  assign T122 = {67'h0, T96};
  assign T96 = T70[1'h0:1'h0];
  assign T97 = 68'h0 - T123;
  assign T123 = {67'h0, T98};
  assign T98 = T70[1'h1:1'h1];
  assign T99 = {T100, T100};
  assign T100 = io_write_bits_data[8'h87:7'h44];
  assign T101 = T103 & T102;
  assign T102 = io_write_bits_wmask[1'h1:1'h1];
  assign T103 = T104 & io_write_valid;
  assign T104 = T70 != 2'h0;
  assign T106 = T107 ? raddr : R105;
  assign io_resp_3 = T109;
  assign T109 = T110;
  assign T110 = {T115, T111};
  assign T111 = T113 ? T115 : T112;
  assign T112 = T62[8'h87:7'h44];
  assign T113 = T114;
  assign T114 = R86[2'h3:2'h3];
  assign T115 = T89[8'h87:7'h44];
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T23) begin
      R21 <= raddr;
    end
    if(io_read_valid) begin
      R28 <= io_read_bits_addr;
    end
    if(T49) begin
      R47 <= raddr;
    end
    if(T81) begin
      R79 <= raddr;
    end
    if(io_read_valid) begin
      R86 <= io_read_bits_addr;
    end
    if(T107) begin
      R105 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input [3:0] io_in_3_bits_way_en,
    input [12:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [3:0] io_in_2_bits_way_en,
    input [12:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [12:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [12:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[12:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[12:0] T2;
  wire[12:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[12:0] T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 2'h0 : T0;
  assign T0 = io_in_1_valid ? 2'h1 : T1;
  assign T1 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T2;
  assign T2 = T8 ? T6 : T3;
  assign T3 = T4 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T4 = T5[1'h0:1'h0];
  assign T5 = chosen;
  assign T6 = T7 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T7 = T5[1'h0:1'h0];
  assign T8 = T5[1'h1:1'h1];
  assign io_out_bits_way_en = T9;
  assign T9 = T14 ? T12 : T10;
  assign T10 = T11 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T11 = T5[1'h0:1'h0];
  assign T12 = T13 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T13 = T5[1'h0:1'h0];
  assign T14 = T5[1'h1:1'h1];
  assign io_out_valid = T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T5[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T5[1'h0:1'h0];
  assign T20 = T5[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T21;
  assign T21 = T22 & io_out_ready;
  assign T22 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 | io_in_2_valid;
  assign T29 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [3:0] io_in_1_bits_way_en,
    input [12:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [135:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [3:0] io_in_0_bits_way_en,
    input [12:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [135:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[3:0] io_out_bits_way_en,
    output[12:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[135:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[135:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[12:0] T3;
  wire[3:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T0;
  assign T0 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T1 = chosen;
  assign io_out_bits_wmask = T2;
  assign T2 = T1 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T3;
  assign T3 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T4;
  assign T4 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [3:0] io_cmd,
    input [3:0] io_typ,
    input [67:0] io_lhs,
    input [67:0] io_rhs,
    output[67:0] io_out
);

  wire[67:0] T125;
  wire[87:0] T0;
  wire[87:0] T1;
  wire[87:0] T126;
  wire[87:0] T2;
  wire[87:0] wmask;
  wire[87:0] T3;
  wire[87:0] T4;
  wire[47:0] T5;
  wire[23:0] T6;
  wire[15:0] T7;
  wire[7:0] T8;
  wire[7:0] T127;
  wire T9;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[10:0] T128;
  wire[8:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[10:0] T129;
  wire[7:0] T25;
  wire[2:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[7:0] T30;
  wire[7:0] T130;
  wire T31;
  wire[7:0] T32;
  wire[7:0] T131;
  wire T33;
  wire[23:0] T34;
  wire[15:0] T35;
  wire[7:0] T36;
  wire[7:0] T132;
  wire T37;
  wire[7:0] T38;
  wire[7:0] T133;
  wire T39;
  wire[7:0] T40;
  wire[7:0] T134;
  wire T41;
  wire[39:0] T42;
  wire[23:0] T43;
  wire[15:0] T44;
  wire[7:0] T45;
  wire[7:0] T135;
  wire T46;
  wire[7:0] T47;
  wire[7:0] T136;
  wire T48;
  wire[7:0] T49;
  wire[7:0] T137;
  wire T50;
  wire[15:0] T51;
  wire[7:0] T52;
  wire[7:0] T138;
  wire T53;
  wire[7:0] T54;
  wire[7:0] T139;
  wire T55;
  wire[87:0] T140;
  wire[67:0] T56;
  wire[3:0] T57;
  wire T58;
  wire[87:0] T59;
  wire[87:0] T141;
  wire[67:0] out;
  wire[67:0] T60;
  wire[67:0] T61;
  wire[67:0] T62;
  wire[67:0] T63;
  wire[67:0] T64;
  wire[67:0] T65;
  wire[67:0] T66;
  wire[67:0] rhs;
  wire[67:0] T142;
  wire[63:0] T67;
  wire[31:0] T68;
  wire[67:0] T143;
  wire[63:0] T69;
  wire[31:0] T70;
  wire[15:0] T71;
  wire[67:0] T144;
  wire[63:0] T72;
  wire[31:0] T73;
  wire[15:0] T74;
  wire[7:0] T75;
  wire[67:0] T76;
  wire[3:0] T77;
  wire T78;
  wire max;
  wire T79;
  wire[4:0] T145;
  wire T80;
  wire[4:0] T146;
  wire min;
  wire T81;
  wire[4:0] T147;
  wire T82;
  wire[4:0] T148;
  wire less;
  wire T83;
  wire cmp_rhs;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire word;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire cmp_lhs;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire sgned;
  wire T100;
  wire[4:0] T149;
  wire T101;
  wire[4:0] T150;
  wire lt;
  wire T102;
  wire T103;
  wire lt_lo;
  wire[31:0] T104;
  wire[31:0] T105;
  wire eq_hi;
  wire[31:0] T106;
  wire[31:0] T107;
  wire lt_hi;
  wire[31:0] T108;
  wire[31:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[67:0] T113;
  wire T114;
  wire[4:0] T151;
  wire[67:0] T115;
  wire T116;
  wire[4:0] T152;
  wire[67:0] T117;
  wire T118;
  wire[4:0] T153;
  wire[67:0] adder_out;
  wire[67:0] T119;
  wire[67:0] T154;
  wire[63:0] mask;
  wire[63:0] T155;
  wire[31:0] T120;
  wire T121;
  wire[3:0] T156;
  wire T157;
  wire[67:0] T122;
  wire[67:0] T123;
  wire[67:0] T158;
  wire[3:0] T159;
  wire T160;
  wire T124;
  wire[4:0] T161;


  assign io_out = T125;
  assign T125 = T0[7'h43:1'h0];
  assign T0 = T59 | T1;
  assign T1 = T2 & T126;
  assign T126 = {20'h0, io_lhs};
  assign T2 = ~ wmask;
  assign wmask = T58 ? T140 : T3;
  assign T3 = T4;
  assign T4 = {T42, T5};
  assign T5 = {T34, T6};
  assign T6 = {T32, T7};
  assign T7 = {T30, T8};
  assign T8 = 8'h0 - T127;
  assign T127 = {7'h0, T9};
  assign T9 = T10[1'h0:1'h0];
  assign T10 = T27 ? T129 : T11;
  assign T11 = T22 ? T128 : T12;
  assign T12 = T16 ? T13 : 11'hff;
  assign T13 = 4'hf << T14;
  assign T14 = {T15, 2'h0};
  assign T15 = io_addr[2'h2:2'h2];
  assign T16 = T18 | T17;
  assign T17 = io_typ == 4'h6;
  assign T18 = io_typ == 4'h2;
  assign T128 = {2'h0, T19};
  assign T19 = 2'h3 << T20;
  assign T20 = {T21, 1'h0};
  assign T21 = io_addr[2'h2:1'h1];
  assign T22 = T24 | T23;
  assign T23 = io_typ == 4'h5;
  assign T24 = io_typ == 4'h1;
  assign T129 = {3'h0, T25};
  assign T25 = 1'h1 << T26;
  assign T26 = io_addr[2'h2:1'h0];
  assign T27 = T29 | T28;
  assign T28 = io_typ == 4'h4;
  assign T29 = io_typ == 4'h0;
  assign T30 = 8'h0 - T130;
  assign T130 = {7'h0, T31};
  assign T31 = T10[1'h1:1'h1];
  assign T32 = 8'h0 - T131;
  assign T131 = {7'h0, T33};
  assign T33 = T10[2'h2:2'h2];
  assign T34 = {T40, T35};
  assign T35 = {T38, T36};
  assign T36 = 8'h0 - T132;
  assign T132 = {7'h0, T37};
  assign T37 = T10[2'h3:2'h3];
  assign T38 = 8'h0 - T133;
  assign T133 = {7'h0, T39};
  assign T39 = T10[3'h4:3'h4];
  assign T40 = 8'h0 - T134;
  assign T134 = {7'h0, T41};
  assign T41 = T10[3'h5:3'h5];
  assign T42 = {T51, T43};
  assign T43 = {T49, T44};
  assign T44 = {T47, T45};
  assign T45 = 8'h0 - T135;
  assign T135 = {7'h0, T46};
  assign T46 = T10[3'h6:3'h6];
  assign T47 = 8'h0 - T136;
  assign T136 = {7'h0, T48};
  assign T48 = T10[3'h7:3'h7];
  assign T49 = 8'h0 - T137;
  assign T137 = {7'h0, T50};
  assign T50 = T10[4'h8:4'h8];
  assign T51 = {T54, T52};
  assign T52 = 8'h0 - T138;
  assign T138 = {7'h0, T53};
  assign T53 = T10[4'h9:4'h9];
  assign T54 = 8'h0 - T139;
  assign T139 = {7'h0, T55};
  assign T55 = T10[4'ha:4'ha];
  assign T140 = {20'h0, T56};
  assign T56 = T57 << 7'h40;
  assign T57 = 4'hf;
  assign T58 = io_typ == 4'hf;
  assign T59 = wmask & T141;
  assign T141 = {20'h0, out};
  assign out = T124 ? adder_out : T60;
  assign T60 = T118 ? T117 : T61;
  assign T61 = T116 ? T115 : T62;
  assign T62 = T114 ? T113 : T63;
  assign T63 = T78 ? io_lhs : T64;
  assign T64 = T58 ? T76 : T65;
  assign T65 = T27 ? T144 : T66;
  assign T66 = T22 ? T143 : rhs;
  assign rhs = T16 ? T142 : io_rhs;
  assign T142 = {4'h0, T67};
  assign T67 = {T68, T68};
  assign T68 = io_rhs[5'h1f:1'h0];
  assign T143 = {4'h0, T69};
  assign T69 = {T70, T70};
  assign T70 = {T71, T71};
  assign T71 = io_rhs[4'hf:1'h0];
  assign T144 = {4'h0, T72};
  assign T72 = {T73, T73};
  assign T73 = {T74, T74};
  assign T74 = {T75, T75};
  assign T75 = io_rhs[3'h7:1'h0];
  assign T76 = T77 << 7'h40;
  assign T77 = io_rhs[2'h3:1'h0];
  assign T78 = less ? min : max;
  assign max = T80 | T79;
  assign T79 = T145 == 5'hf;
  assign T145 = {1'h0, io_cmd};
  assign T80 = T146 == 5'hd;
  assign T146 = {1'h0, io_cmd};
  assign min = T82 | T81;
  assign T81 = T147 == 5'he;
  assign T147 = {1'h0, io_cmd};
  assign T82 = T148 == 5'hc;
  assign T148 = {1'h0, io_cmd};
  assign less = T112 ? lt : T83;
  assign T83 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T86 ? T85 : T84;
  assign T84 = rhs[6'h3f:6'h3f];
  assign T85 = rhs[5'h1f:5'h1f];
  assign T86 = word & T87;
  assign T87 = T88 ^ 1'h1;
  assign T88 = io_addr[2'h2:2'h2];
  assign word = T90 | T89;
  assign T89 = io_typ == 4'h4;
  assign T90 = T92 | T91;
  assign T91 = io_typ == 4'h0;
  assign T92 = T94 | T93;
  assign T93 = io_typ == 4'h6;
  assign T94 = io_typ == 4'h2;
  assign cmp_lhs = T97 ? T96 : T95;
  assign T95 = io_lhs[6'h3f:6'h3f];
  assign T96 = io_lhs[5'h1f:5'h1f];
  assign T97 = word & T98;
  assign T98 = T99 ^ 1'h1;
  assign T99 = io_addr[2'h2:2'h2];
  assign sgned = T101 | T100;
  assign T100 = T149 == 5'hd;
  assign T149 = {1'h0, io_cmd};
  assign T101 = T150 == 5'hc;
  assign T150 = {1'h0, io_cmd};
  assign lt = word ? T110 : T102;
  assign T102 = lt_hi | T103;
  assign T103 = eq_hi & lt_lo;
  assign lt_lo = T105 < T104;
  assign T104 = rhs[5'h1f:1'h0];
  assign T105 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T107 == T106;
  assign T106 = rhs[6'h3f:6'h20];
  assign T107 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T109 < T108;
  assign T108 = rhs[6'h3f:6'h20];
  assign T109 = io_lhs[6'h3f:6'h20];
  assign T110 = T111 ? lt_hi : lt_lo;
  assign T111 = io_addr[2'h2:2'h2];
  assign T112 = cmp_lhs == cmp_rhs;
  assign T113 = io_lhs ^ rhs;
  assign T114 = T151 == 5'h9;
  assign T151 = {1'h0, io_cmd};
  assign T115 = io_lhs | rhs;
  assign T116 = T152 == 5'ha;
  assign T152 = {1'h0, io_cmd};
  assign T117 = io_lhs & rhs;
  assign T118 = T153 == 5'hb;
  assign T153 = {1'h0, io_cmd};
  assign adder_out = T122 + T119;
  assign T119 = rhs & T154;
  assign T154 = {T156, mask};
  assign mask = 64'hffffffffffffffff ^ T155;
  assign T155 = {32'h0, T120};
  assign T120 = T121 << 5'h1f;
  assign T121 = io_addr[2'h2:2'h2];
  assign T156 = T157 ? 4'hf : 4'h0;
  assign T157 = mask[6'h3f:6'h3f];
  assign T122 = T123;
  assign T123 = io_lhs & T158;
  assign T158 = {T159, mask};
  assign T159 = T160 ? 4'hf : 4'h0;
  assign T160 = mask[6'h3f:6'h3f];
  assign T124 = T161 == 5'h8;
  assign T161 = {1'h0, io_cmd};
endmodule

module LockingArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [135:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [135:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[135:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T35;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  locked;
  wire T36;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  reg [1:0] R20;
  wire[1:0] T37;
  wire[1:0] T21;
  wire[2:0] T22;
  wire T23;
  wire[135:0] T24;
  wire[1:0] T25;
  wire[25:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R20 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T35 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T14 & T7;
  assign T7 = T9 | T8;
  assign T8 = 3'h3 == io_out_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h2 == io_out_bits_r_type;
  assign T11 = T13 | T12;
  assign T12 = 3'h1 == io_out_bits_r_type;
  assign T13 = 3'h0 == io_out_bits_r_type;
  assign T14 = io_out_ready & io_out_valid;
  assign T36 = reset ? 1'h0 : T15;
  assign T15 = T17 ? 1'h0 : T16;
  assign T16 = T4 ? 1'h1 : locked;
  assign T17 = T14 & T18;
  assign T18 = T19 == 2'h0;
  assign T19 = R20 + 2'h1;
  assign T37 = reset ? 2'h0 : T21;
  assign T21 = T6 ? T19 : R20;
  assign io_out_bits_r_type = T22;
  assign T22 = T23 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T23 = chosen;
  assign io_out_bits_data = T24;
  assign T24 = T23 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T25;
  assign T25 = T23 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T26;
  assign T26 = T23 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T27;
  assign T27 = T23 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = locked ? T30 : 1'h1;
  assign T30 = lockIdx == 1'h0;
  assign io_in_1_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = locked ? T34 : T33;
  assign T33 = io_in_0_valid ^ 1'h1;
  assign T34 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T17) begin
      locked <= 1'h0;
    end else if(T4) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R20 <= 2'h0;
    end else if(T6) begin
      R20 <= T19;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input  io_cpu_req_bits_kill,
    input [3:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_phys,
    input [43:0] io_cpu_req_bits_addr,
    input [7:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    input [63:0] io_cpu_req_bits_data,
    output io_cpu_resp_valid,
    output[63:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output[3:0] io_cpu_resp_bits_typ,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[7:0] io_cpu_resp_bits_tag,
    output[3:0] io_cpu_resp_bits_cmd,
    output[43:0] io_cpu_resp_bits_addr,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[7:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    output io_cpu_ordered,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[135:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[128:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_header_src,
    output[1:0] io_mem_release_bits_header_dst,
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[135:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[67:0] T564;
  reg [63:0] s2_req_data;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  reg  s1_replay;
  wire T565;
  wire T10;
  wire T11;
  wire s1_write;
  wire T12;
  wire T13;
  reg [4:0] s1_req_cmd;
  wire[4:0] T14;
  wire[4:0] T15;
  wire[4:0] T16;
  reg [4:0] s2_req_cmd;
  wire[4:0] T17;
  wire s2_recycle;
  wire T18;
  reg  s2_recycle_next;
  wire T566;
  wire T19;
  wire T20;
  wire T21;
  reg  s1_valid;
  wire T567;
  wire T22;
  wire T23;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire[1:0] T24;
  wire T25;
  wire s2_hit;
  wire T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  reg [1:0] R40;
  wire[1:0] T41;
  wire T42;
  reg [3:0] s2_tag_match_way;
  wire[3:0] T43;
  wire[3:0] s1_tag_match_way;
  wire[3:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire[3:0] s1_tag_eq_way;
  wire[3:0] T49;
  wire[1:0] T50;
  wire T51;
  wire[18:0] T52;
  wire[31:0] s1_addr;
  wire[12:0] T53;
  reg [43:0] s1_req_addr;
  wire[43:0] T54;
  wire[43:0] T55;
  wire[43:0] T56;
  wire[43:0] T57;
  wire[43:0] T58;
  wire[43:0] T568;
  wire[31:0] T59;
  wire[25:0] T60;
  wire[43:0] T569;
  wire[31:0] T61;
  wire[25:0] T62;
  reg [43:0] s2_req_addr;
  wire[43:0] T63;
  wire[43:0] T570;
  wire T64;
  wire[18:0] T65;
  wire[1:0] T66;
  wire T67;
  wire[18:0] T68;
  wire T69;
  wire[18:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire[1:0] T83;
  reg [1:0] R84;
  wire[1:0] T85;
  wire T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  reg [1:0] R90;
  wire[1:0] T91;
  wire T92;
  wire[1:0] T93;
  wire[1:0] T94;
  reg [1:0] R95;
  wire[1:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire s2_tag_match;
  wire T115;
  wire s2_replay;
  wire T116;
  reg  R117;
  wire T571;
  reg  s2_valid;
  wire T572;
  wire s1_valid_masked;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T123;
  wire[63:0] T124;
  wire[63:0] T125;
  wire T126;
  reg  s1_recycled;
  wire T127;
  wire[67:0] s2_data_word;
  wire[67:0] s2_data_word_prebypass;
  wire[67:0] T128;
  wire[135:0] s2_data_muxed;
  wire[135:0] T129;
  wire[135:0] s2_data_3;
  wire[135:0] T130;
  wire[135:0] T131;
  reg [67:0] R132;
  wire[67:0] T573;
  wire[135:0] T133;
  wire[135:0] T574;
  wire[135:0] T134;
  wire T135;
  wire T136;
  reg [67:0] R137;
  wire[67:0] T138;
  wire[67:0] T139;
  wire T140;
  wire s1_writeback;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[135:0] T145;
  wire[135:0] T146;
  wire[135:0] s2_data_2;
  wire[135:0] T147;
  wire[135:0] T148;
  reg [67:0] R149;
  wire[67:0] T575;
  wire[135:0] T150;
  wire[135:0] T576;
  wire[135:0] T151;
  wire T152;
  wire T153;
  reg [67:0] R154;
  wire[67:0] T155;
  wire[67:0] T156;
  wire T157;
  wire T158;
  wire[135:0] T159;
  wire[135:0] T160;
  wire[135:0] s2_data_1;
  wire[135:0] T161;
  wire[135:0] T162;
  reg [67:0] R163;
  wire[67:0] T577;
  wire[135:0] T164;
  wire[135:0] T578;
  wire[135:0] T165;
  wire T166;
  wire T167;
  reg [67:0] R168;
  wire[67:0] T169;
  wire[67:0] T170;
  wire T171;
  wire T172;
  wire[135:0] T173;
  wire[135:0] s2_data_0;
  wire[135:0] T174;
  wire[135:0] T175;
  reg [67:0] R176;
  wire[67:0] T579;
  wire[135:0] T177;
  wire[135:0] T580;
  wire[135:0] T178;
  wire T179;
  wire T180;
  reg [67:0] R181;
  wire[67:0] T182;
  wire[67:0] T183;
  wire T184;
  wire T185;
  wire[67:0] T186;
  wire T187;
  reg [67:0] s2_store_bypass_data;
  wire[67:0] T188;
  wire[67:0] T189;
  wire[67:0] T190;
  reg [67:0] s4_req_data_;
  wire[67:0] T191;
  wire T192;
  reg  s3_valid;
  wire T581;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire s2_sc_fail;
  wire T203;
  wire s2_lrsc_addr_match;
  wire T204;
  wire[37:0] T205;
  reg [37:0] lrsc_addr;
  wire[37:0] T206;
  wire[37:0] T207;
  wire T208;
  wire s2_lr;
  wire T209;
  wire T210;
  wire s2_valid_masked;
  wire T211;
  wire T212;
  wire s2_nack;
  wire s2_nack_miss;
  wire T213;
  wire T214;
  wire T215;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T216;
  wire s1_nack;
  wire T217;
  wire T218;
  wire T219;
  wire[6:0] T220;
  wire T221;
  wire T222;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T582;
  wire[4:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[4:0] T226;
  wire[4:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire s2_sc;
  wire T231;
  wire T232;
  reg [67:0] s3_req_data_;
  wire[67:0] T233;
  wire[67:0] T234;
  wire[67:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  reg [4:0] s3_req_cmd;
  wire[4:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire[40:0] T258;
  reg [43:0] s3_req_addr;
  wire[43:0] T259;
  wire[40:0] T583;
  wire[28:0] T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire[40:0] T271;
  wire[40:0] T584;
  wire[28:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  reg [4:0] s4_req_cmd;
  wire[4:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire[40:0] T290;
  reg [43:0] s4_req_addr;
  wire[43:0] T291;
  wire[40:0] T585;
  wire[28:0] T292;
  reg  s4_valid;
  wire T586;
  wire T293;
  reg  s2_store_bypass;
  wire T294;
  wire T295;
  reg [3:0] s2_req_typ;
  wire[3:0] T296;
  reg [3:0] s1_req_typ;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[3:0] T587;
  wire[5:0] T588;
  wire[135:0] T300;
  wire[1:0] T301;
  wire T302;
  wire T303;
  wire[12:0] T589;
  reg [3:0] s3_way;
  wire[3:0] T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire[12:0] T590;
  wire[12:0] T591;
  wire[12:0] T592;
  wire[135:0] T312;
  wire[135:0] T313;
  wire[67:0] wdata_encoded_0;
  wire[67:0] wdata_encoded_1;
  wire[6:0] T593;
  wire[37:0] T314;
  wire[6:0] T594;
  wire[37:0] T315;
  reg  s1_req_phys;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  reg  s2_req_phys;
  wire T321;
  wire[30:0] T322;
  wire T323;
  wire T324;
  wire T325;
  wire s1_readwrite;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire s1_read;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire[3:0] T338;
  wire[3:0] s2_replaced_way_en;
  reg [1:0] R339;
  wire[1:0] T340;
  wire[1:0] T341;
  reg [15:0] R342;
  wire[15:0] T595;
  wire[15:0] T343;
  wire[15:0] T344;
  wire[14:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire[1:0] T355;
  wire[1:0] T356;
  wire[20:0] T357;
  wire[20:0] T358;
  wire[20:0] T359;
  wire[20:0] T360;
  reg [1:0] R361;
  wire[1:0] T362;
  wire T363;
  wire T364;
  wire[3:0] s1_replaced_way_en;
  wire[1:0] T365;
  reg [18:0] R366;
  wire[18:0] T367;
  wire T368;
  wire[20:0] T369;
  wire[20:0] T370;
  wire[20:0] T371;
  wire[20:0] T372;
  reg [1:0] R373;
  wire[1:0] T374;
  wire T375;
  wire T376;
  reg [18:0] R377;
  wire[18:0] T378;
  wire T379;
  wire[20:0] T380;
  wire[20:0] T381;
  wire[20:0] T382;
  wire[20:0] T383;
  reg [1:0] R384;
  wire[1:0] T385;
  wire T386;
  wire T387;
  reg [18:0] R388;
  wire[18:0] T389;
  wire T390;
  wire[20:0] T391;
  wire[20:0] T392;
  wire[20:0] T393;
  reg [1:0] R394;
  wire[1:0] T395;
  wire T396;
  wire T397;
  reg [18:0] R398;
  wire[18:0] T399;
  wire T400;
  wire[1:0] T401;
  wire[18:0] T402;
  wire[18:0] T403;
  wire[18:0] T404;
  reg [7:0] s2_req_tag;
  wire[7:0] T405;
  reg [7:0] s1_req_tag;
  wire[7:0] T406;
  wire[7:0] T407;
  wire[7:0] T408;
  reg  s2_req_kill;
  wire T409;
  reg  s1_req_kill;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] probe_bits_p_type;
  wire[25:0] probe_bits_addr;
  wire T436;
  wire T437;
  wire probe_valid;
  wire[135:0] T438;
  wire[135:0] T439;
  wire[2:0] T440;
  wire[135:0] T441;
  wire[1:0] T442;
  wire[25:0] T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire probe_ready;
  wire T447;
  wire T448;
  wire[128:0] T449;
  wire[1:0] T450;
  wire T451;
  wire[135:0] T452;
  wire[1:0] T453;
  wire[25:0] T454;
  wire[1:0] T455;
  wire[1:0] T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire misaligned;
  wire T465;
  wire T466;
  wire[2:0] T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire[1:0] T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire s1_sc;
  wire[3:0] T596;
  wire[63:0] T487;
  wire[63:0] T597;
  wire[63:0] T488;
  wire[63:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[63:0] T493;
  wire[15:0] T494;
  wire[15:0] T495;
  wire[63:0] T496;
  wire[31:0] T497;
  wire[31:0] T498;
  wire[31:0] T499;
  wire T500;
  wire[31:0] T501;
  wire[31:0] T502;
  wire[31:0] T503;
  wire[31:0] T598;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[15:0] T516;
  wire T517;
  wire[47:0] T518;
  wire[47:0] T519;
  wire[47:0] T520;
  wire[47:0] T599;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[7:0] T526;
  wire T527;
  wire[55:0] T528;
  wire[55:0] T529;
  wire[55:0] T530;
  wire[55:0] T600;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire[63:0] T537;
  wire[3:0] T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  reg  block_miss;
  wire T601;
  wire T562;
  wire T563;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[6:0] wb_io_meta_read_bits_idx;
  wire[18:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire[3:0] wb_io_data_req_bits_way_en;
  wire[12:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[25:0] wb_io_release_bits_addr;
  wire[1:0] wb_io_release_bits_client_xact_id;
  wire[135:0] wb_io_release_bits_data;
  wire[2:0] wb_io_release_bits_r_type;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[25:0] prober_io_rep_bits_addr;
  wire[1:0] prober_io_rep_bits_client_xact_id;
  wire[135:0] prober_io_rep_bits_data;
  wire[2:0] prober_io_rep_bits_r_type;
  wire prober_io_meta_read_valid;
  wire[6:0] prober_io_meta_read_bits_idx;
  wire[18:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[6:0] prober_io_meta_write_bits_idx;
  wire[3:0] prober_io_meta_write_bits_way_en;
  wire[18:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[18:0] prober_io_wb_req_bits_tag;
  wire[6:0] prober_io_wb_req_bits_idx;
  wire[3:0] prober_io_wb_req_bits_way_en;
  wire[1:0] prober_io_wb_req_bits_client_xact_id;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[18:0] meta_io_resp_3_tag;
  wire[1:0] meta_io_resp_3_coh_state;
  wire[18:0] meta_io_resp_2_tag;
  wire[1:0] meta_io_resp_2_coh_state;
  wire[18:0] meta_io_resp_1_tag;
  wire[1:0] meta_io_resp_1_coh_state;
  wire[18:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[6:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[6:0] metaWriteArb_io_out_bits_idx;
  wire[3:0] metaWriteArb_io_out_bits_way_en;
  wire[18:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[135:0] data_io_resp_3;
  wire[135:0] data_io_resp_2;
  wire[135:0] data_io_resp_1;
  wire[135:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire[3:0] readArb_io_out_bits_way_en;
  wire[12:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire[3:0] writeArb_io_out_bits_way_en;
  wire[12:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[135:0] writeArb_io_out_bits_data;
  wire[67:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[25:0] releaseArb_io_out_bits_addr;
  wire[1:0] releaseArb_io_out_bits_client_xact_id;
  wire[135:0] releaseArb_io_out_bits_data;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire ser_io_in_ready;
  wire ser_io_out_valid;
  wire[1:0] ser_io_out_bits_header_src;
  wire[1:0] ser_io_out_bits_header_dst;
  wire[135:0] ser_io_out_bits_payload_data;
  wire[1:0] ser_io_out_bits_payload_client_xact_id;
  wire[3:0] ser_io_out_bits_payload_manager_xact_id;
  wire ser_io_out_bits_payload_uncached;
  wire[1:0] ser_io_out_bits_payload_g_type;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[18:0] wbArb_io_out_bits_tag;
  wire[6:0] wbArb_io_out_bits_idx;
  wire[3:0] wbArb_io_out_bits_way_en;
  wire[1:0] wbArb_io_out_bits_client_xact_id;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[18:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[29:0] dtlb_io_ptw_req_bits;
  wire mshrs_io_req_ready;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr;
  wire[1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[135:0] mshrs_io_mem_req_bits_data;
  wire mshrs_io_mem_req_bits_uncached;
  wire[1:0] mshrs_io_mem_req_bits_a_type;
  wire[128:0] mshrs_io_mem_req_bits_subblock;
  wire[3:0] mshrs_io_mem_resp_way_en;
  wire[12:0] mshrs_io_mem_resp_addr;
  wire mshrs_io_meta_read_valid;
  wire[6:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[6:0] mshrs_io_meta_write_bits_idx;
  wire[3:0] mshrs_io_meta_write_bits_way_en;
  wire[18:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire mshrs_io_replay_bits_kill;
  wire[3:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_phys;
  wire[43:0] mshrs_io_replay_bits_addr;
  wire[7:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire[63:0] mshrs_io_replay_bits_data;
  wire mshrs_io_mem_finish_valid;
  wire[1:0] mshrs_io_mem_finish_bits_header_src;
  wire[1:0] mshrs_io_mem_finish_bits_header_dst;
  wire[3:0] mshrs_io_mem_finish_bits_payload_manager_xact_id;
  wire mshrs_io_wb_req_valid;
  wire[18:0] mshrs_io_wb_req_bits_tag;
  wire[6:0] mshrs_io_wb_req_bits_idx;
  wire[3:0] mshrs_io_wb_req_bits_way_en;
  wire[1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    R40 = {1{$random}};
    s2_tag_match_way = {1{$random}};
    s1_req_addr = {2{$random}};
    s2_req_addr = {2{$random}};
    R84 = {1{$random}};
    R90 = {1{$random}};
    R95 = {1{$random}};
    R117 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R132 = {3{$random}};
    R137 = {3{$random}};
    R149 = {3{$random}};
    R154 = {3{$random}};
    R163 = {3{$random}};
    R168 = {3{$random}};
    R176 = {3{$random}};
    R181 = {3{$random}};
    s2_store_bypass_data = {3{$random}};
    s4_req_data_ = {3{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data_ = {3{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R339 = {1{$random}};
    R342 = {1{$random}};
    R361 = {1{$random}};
    R366 = {1{$random}};
    R373 = {1{$random}};
    R377 = {1{$random}};
    R384 = {1{$random}};
    R388 = {1{$random}};
    R394 = {1{$random}};
    R398 = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    block_miss = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = writeArb_io_in_1_ready | T1;
  assign T1 = T2 ^ 1'h1;
  assign T2 = ser_io_out_bits_payload_uncached ? 1'h0 : T3;
  assign T3 = T5 | T4;
  assign T4 = ser_io_out_bits_payload_g_type == 2'h2;
  assign T5 = ser_io_out_bits_payload_g_type == 2'h1;
  assign T6 = io_mem_release_ready;
  assign T564 = {4'h0, s2_req_data};
  assign T7 = T126 ? s1_req_data : T8;
  assign T8 = T11 ? T9 : s2_req_data;
  assign T9 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T565 = reset ? 1'h0 : T10;
  assign T10 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T11 = s1_clk_en & s1_write;
  assign s1_write = T120 | T12;
  assign T12 = T119 | T13;
  assign T13 = s1_req_cmd == 5'h4;
  assign T14 = s2_recycle ? s2_req_cmd : T15;
  assign T15 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T16;
  assign T16 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T17 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T18;
  assign T18 = s2_recycle_ecc | s2_recycle_next;
  assign T566 = reset ? 1'h0 : T19;
  assign T19 = T23 ? T20 : s2_recycle_next;
  assign T20 = T21 & s2_recycle_ecc;
  assign T21 = s1_valid | s1_replay;
  assign T567 = reset ? 1'h0 : T22;
  assign T22 = io_cpu_req_ready & io_cpu_req_valid;
  assign T23 = s1_valid | s1_replay;
  assign s2_recycle_ecc = T25 & s2_data_correctable;
  assign s2_data_correctable = T24[1'h0:1'h0];
  assign T24 = 2'h0;
  assign T25 = T115 & s2_hit;
  assign s2_hit = T98 & T26;
  assign T26 = T36 == T27;
  assign T27 = T28;
  assign T28 = T29 ? 2'h2 : T36;
  assign T29 = T33 | T30;
  assign T30 = T32 | T31;
  assign T31 = s2_req_cmd == 5'h4;
  assign T32 = s2_req_cmd[2'h3:2'h3];
  assign T33 = T35 | T34;
  assign T34 = s2_req_cmd == 5'h7;
  assign T35 = s2_req_cmd == 5'h1;
  assign T36 = T37[1'h1:1'h0];
  assign T37 = T81 | T38;
  assign T38 = T42 ? T39 : 2'h0;
  assign T39 = R40;
  assign T41 = s1_clk_en ? meta_io_resp_3_coh_state : R40;
  assign T42 = s2_tag_match_way[2'h3:2'h3];
  assign T43 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T44;
  assign T44 = {T74, T45};
  assign T45 = {T71, T46};
  assign T46 = T48 & T47;
  assign T47 = meta_io_resp_0_coh_state != 2'h0;
  assign T48 = s1_tag_eq_way[1'h0:1'h0];
  assign s1_tag_eq_way = T49;
  assign T49 = {T66, T50};
  assign T50 = {T64, T51};
  assign T51 = meta_io_resp_0_tag == T52;
  assign T52 = s1_addr >> 4'hd;
  assign s1_addr = {dtlb_io_resp_ppn, T53};
  assign T53 = s1_req_addr[4'hc:1'h0];
  assign T54 = s2_recycle ? s2_req_addr : T55;
  assign T55 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T56;
  assign T56 = prober_io_meta_read_valid ? T569 : T57;
  assign T57 = wb_io_meta_read_valid ? T568 : T58;
  assign T58 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T568 = {12'h0, T59};
  assign T59 = T60 << 3'h6;
  assign T60 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T569 = {12'h0, T61};
  assign T61 = T62 << 3'h6;
  assign T62 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T63 = s1_clk_en ? T570 : s2_req_addr;
  assign T570 = {12'h0, s1_addr};
  assign T64 = meta_io_resp_1_tag == T65;
  assign T65 = s1_addr >> 4'hd;
  assign T66 = {T69, T67};
  assign T67 = meta_io_resp_2_tag == T68;
  assign T68 = s1_addr >> 4'hd;
  assign T69 = meta_io_resp_3_tag == T70;
  assign T70 = s1_addr >> 4'hd;
  assign T71 = T73 & T72;
  assign T72 = meta_io_resp_1_coh_state != 2'h0;
  assign T73 = s1_tag_eq_way[1'h1:1'h1];
  assign T74 = {T78, T75};
  assign T75 = T77 & T76;
  assign T76 = meta_io_resp_2_coh_state != 2'h0;
  assign T77 = s1_tag_eq_way[2'h2:2'h2];
  assign T78 = T80 & T79;
  assign T79 = meta_io_resp_3_coh_state != 2'h0;
  assign T80 = s1_tag_eq_way[2'h3:2'h3];
  assign T81 = T87 | T82;
  assign T82 = T86 ? T83 : 2'h0;
  assign T83 = R84;
  assign T85 = s1_clk_en ? meta_io_resp_2_coh_state : R84;
  assign T86 = s2_tag_match_way[2'h2:2'h2];
  assign T87 = T93 | T88;
  assign T88 = T92 ? T89 : 2'h0;
  assign T89 = R90;
  assign T91 = s1_clk_en ? meta_io_resp_1_coh_state : R90;
  assign T92 = s2_tag_match_way[1'h1:1'h1];
  assign T93 = T97 ? T94 : 2'h0;
  assign T94 = R95;
  assign T96 = s1_clk_en ? meta_io_resp_0_coh_state : R95;
  assign T97 = s2_tag_match_way[1'h0:1'h0];
  assign T98 = s2_tag_match & T99;
  assign T99 = T104 ? T103 : T100;
  assign T100 = T102 | T101;
  assign T101 = T36 == 2'h2;
  assign T102 = T36 == 2'h1;
  assign T103 = T36 == 2'h2;
  assign T104 = T106 | T105;
  assign T105 = s2_req_cmd == 5'h6;
  assign T106 = T108 | T107;
  assign T107 = s2_req_cmd == 5'h3;
  assign T108 = T112 | T109;
  assign T109 = T111 | T110;
  assign T110 = s2_req_cmd == 5'h4;
  assign T111 = s2_req_cmd[2'h3:2'h3];
  assign T112 = T114 | T113;
  assign T113 = s2_req_cmd == 5'h7;
  assign T114 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 4'h0;
  assign T115 = s2_valid | s2_replay;
  assign s2_replay = R117 & T116;
  assign T116 = s2_req_cmd != 5'h5;
  assign T571 = reset ? 1'h0 : s1_replay;
  assign T572 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T118;
  assign T118 = io_cpu_req_bits_kill ^ 1'h1;
  assign T119 = s1_req_cmd[2'h3:2'h3];
  assign T120 = T122 | T121;
  assign T121 = s1_req_cmd == 5'h7;
  assign T122 = s1_req_cmd == 5'h1;
  assign T123 = s2_recycle ? s2_req_data : T124;
  assign T124 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T125;
  assign T125 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T126 = s1_clk_en & s1_recycled;
  assign T127 = s1_clk_en ? s2_recycle : s1_recycled;
  assign s2_data_word = s2_store_bypass ? s2_store_bypass_data : s2_data_word_prebypass;
  assign s2_data_word_prebypass = T187 ? T186 : T128;
  assign T128 = s2_data_muxed[7'h43:1'h0];
  assign s2_data_muxed = T145 | T129;
  assign T129 = T144 ? s2_data_3 : 136'h0;
  assign s2_data_3 = T130;
  assign T130 = T131;
  assign T131 = {R137, R132};
  assign T573 = T133[7'h43:1'h0];
  assign T133 = T135 ? T134 : T574;
  assign T574 = {68'h0, R132};
  assign T134 = data_io_resp_3 >> 1'h0;
  assign T135 = s1_clk_en & T136;
  assign T136 = s1_tag_eq_way[2'h3:2'h3];
  assign T138 = T140 ? T139 : R137;
  assign T139 = data_io_resp_3 >> 7'h44;
  assign T140 = T135 & s1_writeback;
  assign s1_writeback = T142 & T141;
  assign T141 = s1_replay ^ 1'h1;
  assign T142 = s1_clk_en & T143;
  assign T143 = s1_valid ^ 1'h1;
  assign T144 = s2_tag_match_way[2'h3:2'h3];
  assign T145 = T159 | T146;
  assign T146 = T158 ? s2_data_2 : 136'h0;
  assign s2_data_2 = T147;
  assign T147 = T148;
  assign T148 = {R154, R149};
  assign T575 = T150[7'h43:1'h0];
  assign T150 = T152 ? T151 : T576;
  assign T576 = {68'h0, R149};
  assign T151 = data_io_resp_2 >> 1'h0;
  assign T152 = s1_clk_en & T153;
  assign T153 = s1_tag_eq_way[2'h2:2'h2];
  assign T155 = T157 ? T156 : R154;
  assign T156 = data_io_resp_2 >> 7'h44;
  assign T157 = T152 & s1_writeback;
  assign T158 = s2_tag_match_way[2'h2:2'h2];
  assign T159 = T173 | T160;
  assign T160 = T172 ? s2_data_1 : 136'h0;
  assign s2_data_1 = T161;
  assign T161 = T162;
  assign T162 = {R168, R163};
  assign T577 = T164[7'h43:1'h0];
  assign T164 = T166 ? T165 : T578;
  assign T578 = {68'h0, R163};
  assign T165 = data_io_resp_1 >> 1'h0;
  assign T166 = s1_clk_en & T167;
  assign T167 = s1_tag_eq_way[1'h1:1'h1];
  assign T169 = T171 ? T170 : R168;
  assign T170 = data_io_resp_1 >> 7'h44;
  assign T171 = T166 & s1_writeback;
  assign T172 = s2_tag_match_way[1'h1:1'h1];
  assign T173 = T185 ? s2_data_0 : 136'h0;
  assign s2_data_0 = T174;
  assign T174 = T175;
  assign T175 = {R181, R176};
  assign T579 = T177[7'h43:1'h0];
  assign T177 = T179 ? T178 : T580;
  assign T580 = {68'h0, R176};
  assign T178 = data_io_resp_0 >> 1'h0;
  assign T179 = s1_clk_en & T180;
  assign T180 = s1_tag_eq_way[1'h0:1'h0];
  assign T182 = T184 ? T183 : R181;
  assign T183 = data_io_resp_0 >> 7'h44;
  assign T184 = T179 & s1_writeback;
  assign T185 = s2_tag_match_way[1'h0:1'h0];
  assign T186 = s2_data_muxed[8'h87:7'h44];
  assign T187 = 1'h0;
  assign T188 = T276 ? T189 : s2_store_bypass_data;
  assign T189 = T261 ? amoalu_io_out : T190;
  assign T190 = T247 ? s3_req_data_ : s4_req_data_;
  assign T191 = T192 ? s3_req_data_ : s4_req_data_;
  assign T192 = s3_valid & metaReadArb_io_out_valid;
  assign T581 = reset ? 1'h0 : T193;
  assign T193 = T201 & T194;
  assign T194 = T198 | T195;
  assign T195 = T197 | T196;
  assign T196 = s2_req_cmd == 5'h4;
  assign T197 = s2_req_cmd[2'h3:2'h3];
  assign T198 = T200 | T199;
  assign T199 = s2_req_cmd == 5'h7;
  assign T200 = s2_req_cmd == 5'h1;
  assign T201 = T231 & T202;
  assign T202 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T203;
  assign T203 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T204;
  assign T204 = lrsc_addr == T205;
  assign T205 = s2_req_addr >> 3'h6;
  assign T206 = T208 ? T207 : lrsc_addr;
  assign T207 = s2_req_addr >> 3'h6;
  assign T208 = T209 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T209 = T210 | s2_replay;
  assign T210 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T211;
  assign T211 = s2_valid & T212;
  assign T212 = s2_nack ^ 1'h1;
  assign s2_nack = T215 | s2_nack_miss;
  assign s2_nack_miss = T214 & T213;
  assign T213 = mshrs_io_req_ready ^ 1'h1;
  assign T214 = s2_hit ^ 1'h1;
  assign T215 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T216 = T222 ? s1_nack : s2_nack_hit;
  assign s1_nack = T221 | T217;
  assign T217 = T219 & T218;
  assign T218 = prober_io_req_ready ^ 1'h1;
  assign T219 = T220 == prober_io_meta_write_bits_idx;
  assign T220 = s1_req_addr[4'hc:3'h6];
  assign T221 = T323 & dtlb_io_resp_miss;
  assign T222 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T582 = reset ? 5'h0 : T223;
  assign T223 = io_cpu_ptw_sret ? 5'h0 : T224;
  assign T224 = T230 ? 5'h0 : T225;
  assign T225 = T228 ? 5'h1f : T226;
  assign T226 = lrsc_valid ? T227 : lrsc_count;
  assign T227 = lrsc_count - 5'h1;
  assign T228 = T208 & T229;
  assign T229 = lrsc_valid ^ 1'h1;
  assign T230 = T209 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T231 = T232 | s2_replay;
  assign T232 = s2_valid_masked & s2_hit;
  assign T233 = T237 ? T234 : s3_req_data_;
  assign T234 = s2_data_correctable ? T235 : amoalu_io_out;
  assign T235 = T236 ? T186 : T128;
  assign T236 = 1'h0;
  assign T237 = T246 & T238;
  assign T238 = T239 | s2_data_correctable;
  assign T239 = T243 | T240;
  assign T240 = T242 | T241;
  assign T241 = s2_req_cmd == 5'h4;
  assign T242 = s2_req_cmd[2'h3:2'h3];
  assign T243 = T245 | T244;
  assign T244 = s2_req_cmd == 5'h7;
  assign T245 = s2_req_cmd == 5'h1;
  assign T246 = s2_valid | s2_replay;
  assign T247 = T256 & T248;
  assign T248 = T253 | T249;
  assign T249 = T252 | T250;
  assign T250 = s3_req_cmd == 5'h4;
  assign T251 = T237 ? s2_req_cmd : s3_req_cmd;
  assign T252 = s3_req_cmd[2'h3:2'h3];
  assign T253 = T255 | T254;
  assign T254 = s3_req_cmd == 5'h7;
  assign T255 = s3_req_cmd == 5'h1;
  assign T256 = s3_valid & T257;
  assign T257 = T583 == T258;
  assign T258 = s3_req_addr >> 2'h3;
  assign T259 = T237 ? s2_req_addr : s3_req_addr;
  assign T583 = {12'h0, T260};
  assign T260 = s1_addr >> 2'h3;
  assign T261 = T269 & T262;
  assign T262 = T266 | T263;
  assign T263 = T265 | T264;
  assign T264 = s2_req_cmd == 5'h4;
  assign T265 = s2_req_cmd[2'h3:2'h3];
  assign T266 = T268 | T267;
  assign T267 = s2_req_cmd == 5'h7;
  assign T268 = s2_req_cmd == 5'h1;
  assign T269 = T273 & T270;
  assign T270 = T584 == T271;
  assign T271 = s2_req_addr >> 2'h3;
  assign T584 = {12'h0, T272};
  assign T272 = s1_addr >> 2'h3;
  assign T273 = T275 & T274;
  assign T274 = s2_sc_fail ^ 1'h1;
  assign T275 = s2_valid_masked | s2_replay;
  assign T276 = s1_clk_en & T277;
  assign T277 = T293 | T278;
  assign T278 = T288 & T279;
  assign T279 = T285 | T280;
  assign T280 = T284 | T281;
  assign T281 = s4_req_cmd == 5'h4;
  assign T282 = T283 ? s3_req_cmd : s4_req_cmd;
  assign T283 = s3_valid & metaReadArb_io_out_valid;
  assign T284 = s4_req_cmd[2'h3:2'h3];
  assign T285 = T287 | T286;
  assign T286 = s4_req_cmd == 5'h7;
  assign T287 = s4_req_cmd == 5'h1;
  assign T288 = s4_valid & T289;
  assign T289 = T585 == T290;
  assign T290 = s4_req_addr >> 2'h3;
  assign T291 = T283 ? s3_req_addr : s4_req_addr;
  assign T585 = {12'h0, T292};
  assign T292 = s1_addr >> 2'h3;
  assign T586 = reset ? 1'h0 : s3_valid;
  assign T293 = T261 | T247;
  assign T294 = T276 ? 1'h1 : T295;
  assign T295 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T296 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T297 = s2_recycle ? s2_req_typ : T298;
  assign T298 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T299;
  assign T299 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T587 = s2_req_cmd[2'h3:1'h0];
  assign T588 = s2_req_addr[3'h5:1'h0];
  assign T300 = {s3_req_data_, s3_req_data_};
  assign T301 = 1'h1 << T302;
  assign T302 = T303;
  assign T303 = s3_req_addr[2'h3:2'h3];
  assign T589 = s3_req_addr[4'hc:1'h0];
  assign T304 = T237 ? s2_tag_match_way : s3_way;
  assign T305 = ser_io_out_valid & T306;
  assign T306 = ser_io_out_bits_payload_uncached ? 1'h0 : T307;
  assign T307 = T309 | T308;
  assign T308 = ser_io_out_bits_payload_g_type == 2'h2;
  assign T309 = ser_io_out_bits_payload_g_type == 2'h1;
  assign T310 = T311 | T0;
  assign T311 = ser_io_out_valid ^ 1'h1;
  assign T590 = s2_req_addr[4'hc:1'h0];
  assign T591 = mshrs_io_replay_bits_addr[4'hc:1'h0];
  assign T592 = io_cpu_req_bits_addr[4'hc:1'h0];
  assign T312 = T313;
  assign T313 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[7'h43:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[8'h87:7'h44];
  assign T593 = T314[3'h6:1'h0];
  assign T314 = s2_req_addr >> 3'h6;
  assign T594 = T315[3'h6:1'h0];
  assign T315 = io_cpu_req_bits_addr >> 3'h6;
  assign T316 = s2_recycle ? s2_req_phys : T317;
  assign T317 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T318;
  assign T318 = prober_io_meta_read_valid ? 1'h1 : T319;
  assign T319 = wb_io_meta_read_valid ? 1'h1 : T320;
  assign T320 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T321 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T322 = s1_req_addr >> 4'hd;
  assign T323 = T325 & T324;
  assign T324 = s1_req_phys ^ 1'h1;
  assign T325 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T329 | T326;
  assign T326 = T328 | T327;
  assign T327 = s1_req_cmd == 5'h3;
  assign T328 = s1_req_cmd == 5'h2;
  assign T329 = s1_read | s1_write;
  assign s1_read = T333 | T330;
  assign T330 = T332 | T331;
  assign T331 = s1_req_cmd == 5'h4;
  assign T332 = s1_req_cmd[2'h3:2'h3];
  assign T333 = T335 | T334;
  assign T334 = s1_req_cmd == 5'h6;
  assign T335 = s1_req_cmd == 5'h0;
  assign T336 = T0 & ser_io_out_valid;
  assign T337 = io_mem_acquire_ready;
  assign T338 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R339;
  assign T340 = s1_clk_en ? T341 : R339;
  assign T341 = R342[1'h1:1'h0];
  assign T595 = reset ? 16'h1 : T343;
  assign T343 = T353 ? T344 : R342;
  assign T344 = {T346, T345};
  assign T345 = R342[4'hf:1'h1];
  assign T346 = T348 ^ T347;
  assign T347 = R342[3'h5:3'h5];
  assign T348 = T350 ^ T349;
  assign T349 = R342[2'h3:2'h3];
  assign T350 = T352 ^ T351;
  assign T351 = R342[2'h2:2'h2];
  assign T352 = R342[1'h0:1'h0];
  assign T353 = T354;
  assign T354 = mshrs_io_req_ready & T413;
  assign T355 = s2_tag_match ? T401 : T356;
  assign T356 = T357[1'h1:1'h0];
  assign T357 = T369 | T358;
  assign T358 = T368 ? T359 : 21'h0;
  assign T359 = T360;
  assign T360 = {R366, R361};
  assign T362 = T363 ? meta_io_resp_3_coh_state : R361;
  assign T363 = s1_clk_en & T364;
  assign T364 = s1_replaced_way_en[2'h3:2'h3];
  assign s1_replaced_way_en = 1'h1 << T365;
  assign T365 = R342[1'h1:1'h0];
  assign T367 = T363 ? meta_io_resp_3_tag : R366;
  assign T368 = s2_replaced_way_en[2'h3:2'h3];
  assign T369 = T380 | T370;
  assign T370 = T379 ? T371 : 21'h0;
  assign T371 = T372;
  assign T372 = {R377, R373};
  assign T374 = T375 ? meta_io_resp_2_coh_state : R373;
  assign T375 = s1_clk_en & T376;
  assign T376 = s1_replaced_way_en[2'h2:2'h2];
  assign T378 = T375 ? meta_io_resp_2_tag : R377;
  assign T379 = s2_replaced_way_en[2'h2:2'h2];
  assign T380 = T391 | T381;
  assign T381 = T390 ? T382 : 21'h0;
  assign T382 = T383;
  assign T383 = {R388, R384};
  assign T385 = T386 ? meta_io_resp_1_coh_state : R384;
  assign T386 = s1_clk_en & T387;
  assign T387 = s1_replaced_way_en[1'h1:1'h1];
  assign T389 = T386 ? meta_io_resp_1_tag : R388;
  assign T390 = s2_replaced_way_en[1'h1:1'h1];
  assign T391 = T400 ? T392 : 21'h0;
  assign T392 = T393;
  assign T393 = {R398, R394};
  assign T395 = T396 ? meta_io_resp_0_coh_state : R394;
  assign T396 = s1_clk_en & T397;
  assign T397 = s1_replaced_way_en[1'h0:1'h0];
  assign T399 = T396 ? meta_io_resp_0_tag : R398;
  assign T400 = s2_replaced_way_en[1'h0:1'h0];
  assign T401 = T36;
  assign T402 = s2_tag_match ? T404 : T403;
  assign T403 = T357[5'h14:2'h2];
  assign T404 = T403;
  assign T405 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T406 = s2_recycle ? s2_req_tag : T407;
  assign T407 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T408;
  assign T408 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T409 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T410 = s2_recycle ? s2_req_kill : T411;
  assign T411 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T412;
  assign T412 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T413 = s2_nack_hit ? 1'h0 : T414;
  assign T414 = T434 & T415;
  assign T415 = T423 | T416;
  assign T416 = T420 | T417;
  assign T417 = T419 | T418;
  assign T418 = s2_req_cmd == 5'h4;
  assign T419 = s2_req_cmd[2'h3:2'h3];
  assign T420 = T422 | T421;
  assign T421 = s2_req_cmd == 5'h7;
  assign T422 = s2_req_cmd == 5'h1;
  assign T423 = T431 | T424;
  assign T424 = T428 | T425;
  assign T425 = T427 | T426;
  assign T426 = s2_req_cmd == 5'h4;
  assign T427 = s2_req_cmd[2'h3:2'h3];
  assign T428 = T430 | T429;
  assign T429 = s2_req_cmd == 5'h6;
  assign T430 = s2_req_cmd == 5'h0;
  assign T431 = T433 | T432;
  assign T432 = s2_req_cmd == 5'h3;
  assign T433 = s2_req_cmd == 5'h2;
  assign T434 = s2_valid_masked & T435;
  assign T435 = s2_hit ^ 1'h1;
  assign probe_bits_p_type = io_mem_probe_bits_payload_p_type;
  assign probe_bits_addr = io_mem_probe_bits_payload_addr;
  assign T436 = probe_valid & T437;
  assign T437 = lrsc_valid ^ 1'h1;
  assign probe_valid = io_mem_probe_valid;
  assign T438 = T439;
  assign T439 = {T186, T128};
  assign io_mem_release_bits_payload_r_type = T440;
  assign T440 = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_payload_data = T441;
  assign T441 = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_payload_client_xact_id = T442;
  assign T442 = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_payload_addr = T443;
  assign T443 = releaseArb_io_out_bits_addr;
  assign io_mem_release_bits_header_dst = T444;
  assign T444 = 2'h0;
  assign io_mem_release_bits_header_src = T445;
  assign T445 = 2'h0;
  assign io_mem_release_valid = T446;
  assign T446 = releaseArb_io_out_valid;
  assign io_mem_probe_ready = probe_ready;
  assign probe_ready = T447;
  assign T447 = prober_io_req_ready & T448;
  assign T448 = lrsc_valid ^ 1'h1;
  assign io_mem_finish_bits_payload_manager_xact_id = mshrs_io_mem_finish_bits_payload_manager_xact_id;
  assign io_mem_finish_bits_header_dst = mshrs_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = mshrs_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_grant_ready = ser_io_in_ready;
  assign io_mem_acquire_bits_payload_subblock = T449;
  assign T449 = mshrs_io_mem_req_bits_subblock;
  assign io_mem_acquire_bits_payload_a_type = T450;
  assign T450 = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_payload_uncached = T451;
  assign T451 = mshrs_io_mem_req_bits_uncached;
  assign io_mem_acquire_bits_payload_data = T452;
  assign T452 = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_payload_client_xact_id = T453;
  assign T453 = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = T454;
  assign T454 = mshrs_io_mem_req_bits_addr;
  assign io_mem_acquire_bits_header_dst = T455;
  assign T455 = 2'h0;
  assign io_mem_acquire_bits_header_src = T456;
  assign T456 = 2'h0;
  assign io_mem_acquire_valid = T457;
  assign T457 = mshrs_io_mem_req_valid;
  assign io_cpu_ordered = T458;
  assign T458 = T460 & T459;
  assign T459 = s2_valid ^ 1'h1;
  assign T460 = mshrs_io_fence_rdy & T461;
  assign T461 = s1_valid ^ 1'h1;
  assign io_cpu_ptw_req_bits = dtlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_xcpt_pf_st = T462;
  assign T462 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T463;
  assign T463 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T464;
  assign T464 = s1_write & misaligned;
  assign misaligned = T471 | T465;
  assign T465 = T468 & T466;
  assign T466 = T467 != 3'h0;
  assign T467 = s1_req_addr[2'h2:1'h0];
  assign T468 = T470 | T469;
  assign T469 = s1_req_typ == 4'hf;
  assign T470 = s1_req_typ == 4'h3;
  assign T471 = T478 | T472;
  assign T472 = T475 & T473;
  assign T473 = T474 != 2'h0;
  assign T474 = s1_req_addr[1'h1:1'h0];
  assign T475 = T477 | T476;
  assign T476 = s1_req_typ == 4'h6;
  assign T477 = s1_req_typ == 4'h2;
  assign T478 = T481 & T479;
  assign T479 = T480 != 1'h0;
  assign T480 = s1_req_addr[1'h0:1'h0];
  assign T481 = T483 | T482;
  assign T482 = s1_req_typ == 4'h5;
  assign T483 = s1_req_typ == 4'h1;
  assign io_cpu_xcpt_ma_ld = T484;
  assign T484 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T485;
  assign T485 = s1_replay & T486;
  assign T486 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_cmd = T596;
  assign T596 = s2_req_cmd[2'h3:1'h0];
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data_subword = T487;
  assign T487 = T488 | T597;
  assign T597 = {63'h0, s2_sc_fail};
  assign T488 = T539 ? T537 : T489;
  assign T489 = {T528, T490};
  assign T490 = s2_sc ? 8'h0 : T491;
  assign T491 = T527 ? T526 : T492;
  assign T492 = T493[3'h7:1'h0];
  assign T493 = {T518, T494};
  assign T494 = T517 ? T516 : T495;
  assign T495 = T496[4'hf:1'h0];
  assign T496 = {T501, T497};
  assign T497 = T500 ? T499 : T498;
  assign T498 = s2_data_word[5'h1f:1'h0];
  assign T499 = s2_data_word[6'h3f:6'h20];
  assign T500 = s2_req_addr[2'h2:2'h2];
  assign T501 = T513 ? T503 : T502;
  assign T502 = s2_data_word[6'h3f:6'h20];
  assign T503 = 32'h0 - T598;
  assign T598 = {31'h0, T504};
  assign T504 = T506 & T505;
  assign T505 = T497[5'h1f:5'h1f];
  assign T506 = T508 | T507;
  assign T507 = s2_req_typ == 4'h3;
  assign T508 = T510 | T509;
  assign T509 = s2_req_typ == 4'h2;
  assign T510 = T512 | T511;
  assign T511 = s2_req_typ == 4'h1;
  assign T512 = s2_req_typ == 4'h0;
  assign T513 = T515 | T514;
  assign T514 = s2_req_typ == 4'h6;
  assign T515 = s2_req_typ == 4'h2;
  assign T516 = T496[5'h1f:5'h10];
  assign T517 = s2_req_addr[1'h1:1'h1];
  assign T518 = T523 ? T520 : T519;
  assign T519 = T496[6'h3f:5'h10];
  assign T520 = 48'h0 - T599;
  assign T599 = {47'h0, T521};
  assign T521 = T506 & T522;
  assign T522 = T494[4'hf:4'hf];
  assign T523 = T525 | T524;
  assign T524 = s2_req_typ == 4'h5;
  assign T525 = s2_req_typ == 4'h1;
  assign T526 = T493[4'hf:4'h8];
  assign T527 = s2_req_addr[1'h0:1'h0];
  assign T528 = T533 ? T530 : T529;
  assign T529 = T493[6'h3f:4'h8];
  assign T530 = 56'h0 - T600;
  assign T600 = {55'h0, T531};
  assign T531 = T506 & T532;
  assign T532 = T490[3'h7:3'h7];
  assign T533 = s2_sc | T534;
  assign T534 = T536 | T535;
  assign T535 = s2_req_typ == 4'h4;
  assign T536 = s2_req_typ == 4'h0;
  assign T537 = {60'h0, T538};
  assign T538 = s2_data_word[7'h43:7'h40];
  assign T539 = s2_req_typ == 4'hf;
  assign io_cpu_resp_bits_has_data = T540;
  assign T540 = T541 | s2_sc;
  assign T541 = T545 | T542;
  assign T542 = T544 | T543;
  assign T543 = s2_req_cmd == 5'h4;
  assign T544 = s2_req_cmd[2'h3:2'h3];
  assign T545 = T547 | T546;
  assign T546 = s2_req_cmd == 5'h6;
  assign T547 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T548;
  assign T548 = s2_valid & s2_nack;
  assign io_cpu_resp_bits_data = T496;
  assign io_cpu_resp_valid = T549;
  assign T549 = T551 & T550;
  assign T550 = s2_data_correctable ^ 1'h1;
  assign T551 = s2_replay | T552;
  assign T552 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T553;
  assign T553 = block_miss ? 1'h0 : T554;
  assign T554 = T561 ? 1'h0 : T555;
  assign T555 = T560 ? 1'h0 : T556;
  assign T556 = T557 == 1'h0;
  assign T557 = T559 & T558;
  assign T558 = io_cpu_req_bits_phys ^ 1'h1;
  assign T559 = dtlb_io_req_ready ^ 1'h1;
  assign T560 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T561 = readArb_io_in_3_ready ^ 1'h1;
  assign T601 = reset ? 1'h0 : T562;
  assign T562 = T563 & s2_nack_miss;
  assign T563 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_tag( wbArb_io_out_bits_tag ),
       .io_req_bits_idx( wbArb_io_out_bits_idx ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( T438 ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr( wb_io_release_bits_addr ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T436 ),
       .io_req_bits_addr( probe_bits_addr ),
       .io_req_bits_p_type( probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr( prober_io_rep_bits_addr ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_tag( prober_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( prober_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_line_state_state( T36 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign prober.io_req_bits_client_xact_id = {1{$random}};
// synthesis translate_on
`endif
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T413 ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T402 ),
       .io_req_bits_old_meta_coh_state( T355 ),
       .io_req_bits_way_en( T338 ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( T337 ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr( mshrs_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_uncached( mshrs_io_mem_req_bits_uncached ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_subblock( mshrs_io_mem_req_bits_subblock ),
       .io_mem_resp_way_en( mshrs_io_mem_resp_way_en ),
       .io_mem_resp_addr( mshrs_io_mem_resp_addr ),
       //.io_mem_resp_wmask(  )
       //.io_mem_resp_data(  )
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_mem_grant_valid( T336 ),
       .io_mem_grant_bits_header_src( ser_io_out_bits_header_src ),
       .io_mem_grant_bits_header_dst( ser_io_out_bits_header_dst ),
       .io_mem_grant_bits_payload_data( ser_io_out_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( ser_io_out_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( ser_io_out_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( ser_io_out_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( ser_io_out_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( mshrs_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( mshrs_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( mshrs_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( mshrs_io_mem_finish_bits_payload_manager_xact_id ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T323 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T322 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_resp_miss( dtlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits( dtlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_3_tag( meta_io_resp_3_tag ),
       .io_resp_3_coh_state( meta_io_resp_3_coh_state ),
       .io_resp_2_tag( meta_io_resp_2_tag ),
       .io_resp_2_coh_state( meta_io_resp_2_coh_state ),
       .io_resp_1_tag( meta_io_resp_1_tag ),
       .io_resp_1_coh_state( meta_io_resp_1_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T594 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T593 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T312 ),
       .io_resp_3( data_io_resp_3 ),
       .io_resp_2( data_io_resp_2 ),
       .io_resp_1( data_io_resp_1 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 4'hf ),
       .io_in_3_bits_addr( T592 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 4'hf ),
       .io_in_1_bits_addr( T591 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 4'hf ),
       .io_in_0_bits_addr( T590 ),
       .io_out_ready( T310 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T305 ),
       .io_in_1_bits_way_en( mshrs_io_mem_resp_way_en ),
       .io_in_1_bits_addr( mshrs_io_mem_resp_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( ser_io_out_bits_payload_data ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T589 ),
       .io_in_0_bits_wmask( T301 ),
       .io_in_0_bits_data( T300 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T588 ),
       .io_cmd( T587 ),
       .io_typ( s2_req_typ ),
       .io_lhs( s2_data_word ),
       .io_rhs( T564 ),
       .io_out( amoalu_io_out )
  );
  LockingArbiter_0 releaseArb(.clk(clk), .reset(reset),
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr( prober_io_rep_bits_addr ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr( wb_io_release_bits_addr ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_out_ready( T6 ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr( releaseArb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  FlowThroughSerializer ser(
       .io_in_ready( ser_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_manager_xact_id( io_mem_grant_bits_payload_manager_xact_id ),
       .io_in_bits_payload_uncached( io_mem_grant_bits_payload_uncached ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( T0 ),
       .io_out_valid( ser_io_out_valid ),
       .io_out_bits_header_src( ser_io_out_bits_header_src ),
       .io_out_bits_header_dst( ser_io_out_bits_header_dst ),
       .io_out_bits_payload_data( ser_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( ser_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( ser_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( ser_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( ser_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_tag( prober_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( prober_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_tag( wbArb_io_out_bits_tag ),
       .io_out_bits_idx( wbArb_io_out_bits_idx ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(T126) begin
      s2_req_data <= s1_req_data;
    end else if(T11) begin
      s2_req_data <= T9;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T10;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T23) begin
      s2_recycle_next <= T20;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T22;
    end
    if(s1_clk_en) begin
      R40 <= meta_io_resp_3_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T569;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T568;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T570;
    end
    if(s1_clk_en) begin
      R84 <= meta_io_resp_2_coh_state;
    end
    if(s1_clk_en) begin
      R90 <= meta_io_resp_1_coh_state;
    end
    if(s1_clk_en) begin
      R95 <= meta_io_resp_0_coh_state;
    end
    if(reset) begin
      R117 <= 1'h0;
    end else begin
      R117 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R132 <= T573;
    if(T140) begin
      R137 <= T139;
    end
    R149 <= T575;
    if(T157) begin
      R154 <= T156;
    end
    R163 <= T577;
    if(T171) begin
      R168 <= T170;
    end
    R176 <= T579;
    if(T184) begin
      R181 <= T183;
    end
    if(T276) begin
      s2_store_bypass_data <= T189;
    end
    if(T192) begin
      s4_req_data_ <= s3_req_data_;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T193;
    end
    if(T208) begin
      lrsc_addr <= T207;
    end
    if(T222) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_ptw_sret) begin
      lrsc_count <= 5'h0;
    end else if(T230) begin
      lrsc_count <= 5'h0;
    end else if(T228) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T227;
    end
    if(T237) begin
      s3_req_data_ <= T234;
    end
    if(T237) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T237) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T283) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T283) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T276) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T237) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R339 <= T341;
    end
    if(reset) begin
      R342 <= 16'h1;
    end else if(T353) begin
      R342 <= T344;
    end
    if(T363) begin
      R361 <= meta_io_resp_3_coh_state;
    end
    if(T363) begin
      R366 <= meta_io_resp_3_tag;
    end
    if(T375) begin
      R373 <= meta_io_resp_2_coh_state;
    end
    if(T375) begin
      R377 <= meta_io_resp_2_tag;
    end
    if(T386) begin
      R384 <= meta_io_resp_1_coh_state;
    end
    if(T386) begin
      R388 <= meta_io_resp_1_tag;
    end
    if(T396) begin
      R394 <= meta_io_resp_0_coh_state;
    end
    if(T396) begin
      R398 <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T562;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [29:0] io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [29:0] io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output[29:0] io_out_bits,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T25;
  wire T3;
  wire T4;
  wire[29:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T25 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits = T5;
  assign T5 = T6 ? io_in_1_bits : io_in_0_bits;
  assign T6 = chosen;
  assign io_out_valid = T7;
  assign T7 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = T16 | T10;
  assign T10 = T11 ^ 1'h1;
  assign T11 = T14 | T12;
  assign T12 = io_in_1_valid & T13;
  assign T13 = last_grant < 1'h1;
  assign T14 = io_in_0_valid & T15;
  assign T15 = last_grant < 1'h0;
  assign T16 = last_grant < 1'h0;
  assign io_in_1_ready = T17;
  assign T17 = T18 & io_out_ready;
  assign T18 = T22 | T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T21 | io_in_0_valid;
  assign T21 = T14 | T12;
  assign T22 = T24 & T23;
  assign T23 = last_grant < 1'h1;
  assign T24 = T14 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [29:0] io_requestor_1_req_bits,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[18:0] io_requestor_1_resp_bits_ppn,
    output[5:0] io_requestor_1_resp_bits_perm,
    output[7:0] io_requestor_1_status_ip,
    output[7:0] io_requestor_1_status_im,
    output[6:0] io_requestor_1_status_zero,
    output io_requestor_1_status_er,
    output io_requestor_1_status_vm,
    output io_requestor_1_status_s64,
    output io_requestor_1_status_u64,
    output io_requestor_1_status_ef,
    output io_requestor_1_status_pei,
    output io_requestor_1_status_ei,
    output io_requestor_1_status_ps,
    output io_requestor_1_status_s,
    output io_requestor_1_invalidate,
    output io_requestor_1_sret,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [29:0] io_requestor_0_req_bits,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[18:0] io_requestor_0_resp_bits_ppn,
    output[5:0] io_requestor_0_resp_bits_perm,
    output[7:0] io_requestor_0_status_ip,
    output[7:0] io_requestor_0_status_im,
    output[6:0] io_requestor_0_status_zero,
    output io_requestor_0_status_er,
    output io_requestor_0_status_vm,
    output io_requestor_0_status_s64,
    output io_requestor_0_status_u64,
    output io_requestor_0_status_ef,
    output io_requestor_0_status_pei,
    output io_requestor_0_status_ei,
    output io_requestor_0_status_ps,
    output io_requestor_0_status_s,
    output io_requestor_0_invalidate,
    output io_requestor_0_sret,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[3:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    //output[7:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    //output[63:0] io_mem_req_bits_data
    input  io_mem_resp_valid,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [3:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    //input  io_mem_ptw_req_valid
    //input [29:0] io_mem_ptw_req_bits
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_sret,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T75;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  reg [1:0] count;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[43:0] T76;
  wire[31:0] T30;
  wire[28:0] T31;
  wire[28:0] T32;
  wire[9:0] vpn_idx;
  wire[9:0] T33;
  wire[9:0] T34;
  wire[9:0] T35;
  reg [29:0] r_req_vpn;
  wire[29:0] T36;
  wire T37;
  wire[9:0] T38;
  wire[19:0] T39;
  wire T40;
  wire[1:0] T41;
  wire[9:0] T42;
  wire[29:0] T43;
  wire T44;
  wire[18:0] T45;
  reg [63:0] r_pte;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T77;
  wire[31:0] T48;
  wire[12:0] T49;
  wire[18:0] T50;
  wire T51;
  wire[5:0] T52;
  wire[18:0] T78;
  wire[30:0] T53;
  wire[30:0] resp_ppn;
  wire[30:0] T54;
  wire[30:0] T55;
  wire[19:0] T56;
  wire[10:0] T57;
  wire[30:0] T58;
  wire[9:0] T59;
  wire[20:0] T60;
  wire T61;
  wire[1:0] T62;
  wire[30:0] r_resp_ppn;
  wire T63;
  wire resp_err;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  reg  r_req_dest;
  wire T68;
  wire resp_val;
  wire T69;
  wire T70;
  wire[5:0] T71;
  wire[18:0] T79;
  wire[30:0] T72;
  wire T73;
  wire T74;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[29:0] arb_io_out_bits;
  wire arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    r_req_vpn = {1{$random}};
    r_pte = {2{$random}};
    r_req_dest = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = state == 3'h0;
  assign T75 = reset ? 3'h0 : T1;
  assign T1 = T29 ? 3'h0 : T2;
  assign T2 = T28 ? 3'h0 : T3;
  assign T3 = T21 ? 3'h1 : T4;
  assign T4 = T16 ? 3'h3 : T5;
  assign T5 = T15 ? 3'h4 : T6;
  assign T6 = T13 ? 3'h1 : T7;
  assign T7 = T11 ? 3'h2 : T8;
  assign T8 = T9 ? 3'h1 : state;
  assign T9 = T10 & arb_io_out_valid;
  assign T10 = 3'h0 == state;
  assign T11 = T12 & io_mem_req_ready;
  assign T12 = 3'h1 == state;
  assign T13 = T14 & io_mem_resp_bits_nack;
  assign T14 = 3'h2 == state;
  assign T15 = T14 & io_mem_resp_valid;
  assign T16 = T19 & T17;
  assign T17 = T18 ^ 1'h1;
  assign T18 = io_mem_resp_bits_data[1'h1:1'h1];
  assign T19 = T15 & T20;
  assign T20 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T21 = T19 & T22;
  assign T22 = T27 & T23;
  assign T23 = count < 2'h2;
  assign T24 = T21 ? T26 : T25;
  assign T25 = T10 ? 2'h0 : count;
  assign T26 = count + 2'h1;
  assign T27 = T17 ^ 1'h1;
  assign T28 = 3'h3 == state;
  assign T29 = 3'h4 == state;
//  assign io_mem_ptw_sret = {1{$random}};
//  assign io_mem_ptw_invalidate = {1{$random}};
//  assign io_mem_ptw_status_s = {1{$random}};
//  assign io_mem_ptw_status_ps = {1{$random}};
//  assign io_mem_ptw_status_ei = {1{$random}};
//  assign io_mem_ptw_status_pei = {1{$random}};
//  assign io_mem_ptw_status_ef = {1{$random}};
//  assign io_mem_ptw_status_u64 = {1{$random}};
//  assign io_mem_ptw_status_s64 = {1{$random}};
//  assign io_mem_ptw_status_vm = {1{$random}};
//  assign io_mem_ptw_status_er = {1{$random}};
//  assign io_mem_ptw_status_zero = {1{$random}};
//  assign io_mem_ptw_status_im = {1{$random}};
//  assign io_mem_ptw_status_ip = {1{$random}};
//  assign io_mem_ptw_resp_bits_perm = {1{$random}};
//  assign io_mem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_mem_ptw_resp_bits_error = {1{$random}};
//  assign io_mem_ptw_resp_valid = {1{$random}};
//  assign io_mem_ptw_req_ready = {1{$random}};
//  assign io_mem_req_bits_data = {2{$random}};
  assign io_mem_req_bits_cmd = 5'h0;
//  assign io_mem_req_bits_tag = {1{$random}};
  assign io_mem_req_bits_addr = T76;
  assign T76 = {12'h0, T30};
  assign T30 = T31 << 2'h3;
  assign T31 = T32;
  assign T32 = {T45, vpn_idx};
  assign vpn_idx = T44 ? T42 : T33;
  assign T33 = T40 ? T38 : T34;
  assign T34 = T35[4'h9:1'h0];
  assign T35 = r_req_vpn >> 5'h14;
  assign T36 = T37 ? arb_io_out_bits : r_req_vpn;
  assign T37 = T0 & arb_io_out_valid;
  assign T38 = T39[4'h9:1'h0];
  assign T39 = r_req_vpn >> 4'ha;
  assign T40 = T41[1'h0:1'h0];
  assign T41 = count;
  assign T42 = T43[4'h9:1'h0];
  assign T43 = r_req_vpn >> 1'h0;
  assign T44 = T41[1'h1:1'h1];
  assign T45 = r_pte[5'h1f:4'hd];
  assign T46 = io_mem_resp_valid ? io_mem_resp_bits_data : T47;
  assign T47 = T37 ? T77 : r_pte;
  assign T77 = {32'h0, T48};
  assign T48 = {T50, T49};
  assign T49 = io_mem_resp_bits_data[4'hc:1'h0];
  assign T50 = io_dpath_ptbr[5'h1f:4'hd];
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 4'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T51;
  assign T51 = state == 3'h1;
  assign io_requestor_0_sret = io_dpath_sret;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_s = io_dpath_status_s;
  assign io_requestor_0_status_ps = io_dpath_status_ps;
  assign io_requestor_0_status_ei = io_dpath_status_ei;
  assign io_requestor_0_status_pei = io_dpath_status_pei;
  assign io_requestor_0_status_ef = io_dpath_status_ef;
  assign io_requestor_0_status_u64 = io_dpath_status_u64;
  assign io_requestor_0_status_s64 = io_dpath_status_s64;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_er = io_dpath_status_er;
  assign io_requestor_0_status_zero = io_dpath_status_zero;
  assign io_requestor_0_status_im = io_dpath_status_im;
  assign io_requestor_0_status_ip = io_dpath_status_ip;
  assign io_requestor_0_resp_bits_perm = T52;
  assign T52 = r_pte[4'h8:2'h3];
  assign io_requestor_0_resp_bits_ppn = T78;
  assign T78 = T53[5'h12:1'h0];
  assign T53 = resp_ppn;
  assign resp_ppn = T63 ? r_resp_ppn : T54;
  assign T54 = T61 ? T58 : T55;
  assign T55 = {T57, T56};
  assign T56 = r_req_vpn[5'h13:1'h0];
  assign T57 = r_resp_ppn >> 5'h14;
  assign T58 = {T60, T59};
  assign T59 = r_req_vpn[4'h9:1'h0];
  assign T60 = r_resp_ppn >> 4'ha;
  assign T61 = T62[1'h0:1'h0];
  assign T62 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hd;
  assign T63 = T62[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = T65 | T64;
  assign T64 = state == 3'h2;
  assign T65 = state == 3'h4;
  assign io_requestor_0_resp_valid = T66;
  assign T66 = resp_val & T67;
  assign T67 = r_req_dest == 1'h0;
  assign T68 = T37 ? arb_io_chosen : r_req_dest;
  assign resp_val = T70 | T69;
  assign T69 = state == 3'h4;
  assign T70 = state == 3'h3;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_sret = io_dpath_sret;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_s = io_dpath_status_s;
  assign io_requestor_1_status_ps = io_dpath_status_ps;
  assign io_requestor_1_status_ei = io_dpath_status_ei;
  assign io_requestor_1_status_pei = io_dpath_status_pei;
  assign io_requestor_1_status_ef = io_dpath_status_ef;
  assign io_requestor_1_status_u64 = io_dpath_status_u64;
  assign io_requestor_1_status_s64 = io_dpath_status_s64;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_er = io_dpath_status_er;
  assign io_requestor_1_status_zero = io_dpath_status_zero;
  assign io_requestor_1_status_im = io_dpath_status_im;
  assign io_requestor_1_status_ip = io_dpath_status_ip;
  assign io_requestor_1_resp_bits_perm = T71;
  assign T71 = r_pte[4'h8:2'h3];
  assign io_requestor_1_resp_bits_ppn = T79;
  assign T79 = T72[5'h12:1'h0];
  assign T72 = resp_ppn;
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T73;
  assign T73 = resp_val & T74;
  assign T74 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits( io_requestor_1_req_bits ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits( io_requestor_0_req_bits ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits( arb_io_out_bits ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T29) begin
      state <= 3'h0;
    end else if(T28) begin
      state <= 3'h0;
    end else if(T21) begin
      state <= 3'h1;
    end else if(T16) begin
      state <= 3'h3;
    end else if(T15) begin
      state <= 3'h4;
    end else if(T13) begin
      state <= 3'h1;
    end else if(T11) begin
      state <= 3'h2;
    end else if(T9) begin
      state <= 3'h1;
    end
    if(T21) begin
      count <= T26;
    end else if(T10) begin
      count <= 2'h0;
    end
    if(T37) begin
      r_req_vpn <= arb_io_out_bits;
    end
    if(io_mem_resp_valid) begin
      r_pte <= io_mem_resp_bits_data;
    end else if(T37) begin
      r_pte <= T77;
    end
    if(T37) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module Control(input clk, input reset,
    output[2:0] io_dpath_sel_pc,
    output io_dpath_killd,
    output io_dpath_killm,
    output io_dpath_ren_1,
    output io_dpath_ren_0,
    output io_dpath_ex_ctrl_legal,
    output io_dpath_ex_ctrl_fp,
    output io_dpath_ex_ctrl_rocc,
    output io_dpath_ex_ctrl_branch,
    output io_dpath_ex_ctrl_jal,
    output io_dpath_ex_ctrl_jalr,
    output io_dpath_ex_ctrl_rxs2,
    output io_dpath_ex_ctrl_rxs1,
    output[1:0] io_dpath_ex_ctrl_sel_alu2,
    output[1:0] io_dpath_ex_ctrl_sel_alu1,
    output[2:0] io_dpath_ex_ctrl_sel_imm,
    output io_dpath_ex_ctrl_alu_dw,
    output[3:0] io_dpath_ex_ctrl_alu_fn,
    output io_dpath_ex_ctrl_mem,
    output[4:0] io_dpath_ex_ctrl_mem_cmd,
    output[3:0] io_dpath_ex_ctrl_mem_type,
    output io_dpath_ex_ctrl_rfs1,
    output io_dpath_ex_ctrl_rfs2,
    output io_dpath_ex_ctrl_rfs3,
    output io_dpath_ex_ctrl_wfd,
    output io_dpath_ex_ctrl_div,
    output io_dpath_ex_ctrl_wxd,
    output[1:0] io_dpath_ex_ctrl_csr,
    output io_dpath_ex_ctrl_fence_i,
    output io_dpath_ex_ctrl_sret,
    output io_dpath_ex_ctrl_scall,
    output io_dpath_ex_ctrl_fence,
    output io_dpath_ex_ctrl_amo,
    output io_dpath_mem_ctrl_legal,
    output io_dpath_mem_ctrl_fp,
    output io_dpath_mem_ctrl_rocc,
    output io_dpath_mem_ctrl_branch,
    output io_dpath_mem_ctrl_jal,
    output io_dpath_mem_ctrl_jalr,
    output io_dpath_mem_ctrl_rxs2,
    output io_dpath_mem_ctrl_rxs1,
    output[1:0] io_dpath_mem_ctrl_sel_alu2,
    output[1:0] io_dpath_mem_ctrl_sel_alu1,
    output[2:0] io_dpath_mem_ctrl_sel_imm,
    output io_dpath_mem_ctrl_alu_dw,
    output[3:0] io_dpath_mem_ctrl_alu_fn,
    output io_dpath_mem_ctrl_mem,
    output[4:0] io_dpath_mem_ctrl_mem_cmd,
    output[3:0] io_dpath_mem_ctrl_mem_type,
    output io_dpath_mem_ctrl_rfs1,
    output io_dpath_mem_ctrl_rfs2,
    output io_dpath_mem_ctrl_rfs3,
    output io_dpath_mem_ctrl_wfd,
    output io_dpath_mem_ctrl_div,
    output io_dpath_mem_ctrl_wxd,
    output[1:0] io_dpath_mem_ctrl_csr,
    output io_dpath_mem_ctrl_fence_i,
    output io_dpath_mem_ctrl_sret,
    output io_dpath_mem_ctrl_scall,
    output io_dpath_mem_ctrl_fence,
    output io_dpath_mem_ctrl_amo,
    output[2:0] io_dpath_csr,
    output io_dpath_sret,
    output io_dpath_ex_valid,
    output io_dpath_wb_wen,
    output io_dpath_bypass_1,
    output io_dpath_bypass_0,
    output[1:0] io_dpath_bypass_src_1,
    output[1:0] io_dpath_bypass_src_0,
    output io_dpath_ll_ready,
    output io_dpath_retire,
    output io_dpath_exception,
    output[63:0] io_dpath_cause,
    output io_dpath_badvaddr_wen,
    input [31:0] io_dpath_inst,
    input  io_dpath_mem_br_taken,
    input  io_dpath_mem_misprediction,
    input  io_dpath_div_mul_rdy,
    input  io_dpath_ll_wen,
    input [4:0] io_dpath_ll_waddr,
    input [4:0] io_dpath_ex_waddr,
    input  io_dpath_mem_rs1_ra,
    input [4:0] io_dpath_mem_waddr,
    input [4:0] io_dpath_wb_waddr,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s,
    input  io_dpath_fp_sboard_clr,
    input [4:0] io_dpath_fp_sboard_clra,
    input  io_dpath_csr_replay,
    output io_imem_req_valid,
    //output[43:0] io_imem_req_bits_pc
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_btb_update_bits_pc
    //output[42:0] io_imem_btb_update_bits_target
    //output io_imem_btb_update_bits_taken
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    //output[42:0] io_imem_btb_update_bits_br_pc
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output[42:0] io_imem_bht_update_bits_prediction_bits_target,
    output[5:0] io_imem_bht_update_bits_prediction_bits_entry,
    output[6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_bht_update_bits_pc
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    //output[42:0] io_imem_ras_update_bits_returnAddr
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output[42:0] io_imem_ras_update_bits_prediction_bits_target,
    output[5:0] io_imem_ras_update_bits_prediction_bits_entry,
    output[6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[3:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    //output[43:0] io_dmem_req_bits_addr
    //output[7:0] io_dmem_req_bits_tag
    output[4:0] io_dmem_req_bits_cmd,
    //output[63:0] io_dmem_req_bits_data
    input  io_dmem_resp_valid,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [3:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output io_fpu_valid,
    input  io_fpu_fcsr_rdy,
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    input [4:0] io_fpu_dec_cmd,
    input  io_fpu_dec_ldst,
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    input  io_fpu_dec_swap23,
    input  io_fpu_dec_single,
    input  io_fpu_dec_fromint,
    input  io_fpu_dec_toint,
    input  io_fpu_dec_fastpipe,
    input  io_fpu_dec_fma,
    input  io_fpu_dec_round,
    input  io_fpu_sboard_set,
    input  io_fpu_sboard_clr,
    input [4:0] io_fpu_sboard_clra,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [3:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[3:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[135:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_manager_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_manager_xact_id,
    //output io_rocc_dmem_acquire_ready
    input  io_rocc_dmem_acquire_valid,
    input [1:0] io_rocc_dmem_acquire_bits_header_src,
    input [1:0] io_rocc_dmem_acquire_bits_header_dst,
    input [25:0] io_rocc_dmem_acquire_bits_payload_addr,
    input [1:0] io_rocc_dmem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_acquire_bits_payload_data,
    input  io_rocc_dmem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_dmem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_dmem_acquire_bits_payload_subblock,
    input  io_rocc_dmem_grant_ready,
    //output io_rocc_dmem_grant_valid
    //output[1:0] io_rocc_dmem_grant_bits_header_src
    //output[1:0] io_rocc_dmem_grant_bits_header_dst
    //output[135:0] io_rocc_dmem_grant_bits_payload_data
    //output[1:0] io_rocc_dmem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_dmem_grant_bits_payload_manager_xact_id
    //output io_rocc_dmem_grant_bits_payload_uncached
    //output[1:0] io_rocc_dmem_grant_bits_payload_g_type
    //output io_rocc_dmem_finish_ready
    input  io_rocc_dmem_finish_valid,
    input [1:0] io_rocc_dmem_finish_bits_header_src,
    input [1:0] io_rocc_dmem_finish_bits_header_dst,
    input [3:0] io_rocc_dmem_finish_bits_payload_manager_xact_id,
    input  io_rocc_dmem_probe_ready,
    //output io_rocc_dmem_probe_valid
    //output[1:0] io_rocc_dmem_probe_bits_header_src
    //output[1:0] io_rocc_dmem_probe_bits_header_dst
    //output[25:0] io_rocc_dmem_probe_bits_payload_addr
    //output[1:0] io_rocc_dmem_probe_bits_payload_p_type
    //output io_rocc_dmem_release_ready
    input  io_rocc_dmem_release_valid,
    input [1:0] io_rocc_dmem_release_bits_header_src,
    input [1:0] io_rocc_dmem_release_bits_header_dst,
    input [25:0] io_rocc_dmem_release_bits_payload_addr,
    input [1:0] io_rocc_dmem_release_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_release_bits_payload_data,
    input [2:0] io_rocc_dmem_release_bits_payload_r_type,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire T0;
  reg  wb_reg_xcpt;
  wire T1;
  wire T2;
  wire take_pc_wb;
  wire T3;
  wire T4;
  wire replay_wb;
  wire T5;
  wire T6;
  wire T7;
  reg  wb_ctrl_rocc;
  wire T8;
  reg  mem_ctrl_rocc;
  wire T9;
  reg  ex_ctrl_rocc;
  wire T10;
  wire id_ctrl_rocc;
  wire T11;
  wire ctrl_killd;
  wire T12;
  wire ctrl_draind;
  wire id_interrupt_unmasked;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire ctrl_stalld;
  wire id_do_fence;
  wire T44;
  wire id_csr_flush;
  wire T45;
  wire T46;
  wire T47;
  wire[11:0] T48;
  wire[11:0] id_csr_addr;
  wire T49;
  wire[11:0] T50;
  wire T51;
  wire id_csr_wen;
  wire T52;
  wire T53;
  wire T54;
  wire[1:0] id_ctrl_csr;
  wire[1:0] T55;
  wire T56;
  wire[31:0] T57;
  wire T58;
  wire[31:0] T59;
  wire T60;
  wire T61;
  wire[4:0] id_raddr1;
  wire id_csr_en;
  wire T62;
  wire T63;
  wire T64;
  wire id_ctrl_mem;
  wire T65;
  wire T66;
  wire[31:0] T67;
  wire T68;
  wire T69;
  wire[31:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T76;
  wire T77;
  wire T78;
  wire[31:0] T79;
  wire T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire[31:0] T87;
  reg  id_reg_fence;
  wire T905;
  wire T88;
  wire T89;
  wire id_fence_next;
  wire T90;
  wire id_amo_rl;
  wire id_ctrl_amo;
  wire T91;
  wire[31:0] T92;
  wire id_ctrl_fence;
  wire T93;
  wire[31:0] T94;
  wire T95;
  wire id_ctrl_fence_i;
  wire T96;
  wire[31:0] T97;
  wire T98;
  wire id_amo_aq;
  wire id_mem_busy;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire id_stall_fpu;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[4:0] T109;
  wire[4:0] T110;
  wire[4:0] id_waddr;
  wire T111;
  reg [31:0] R112;
  wire[31:0] T906;
  wire[31:0] T113;
  wire[31:0] T114;
  wire[31:0] T115;
  wire[31:0] T116;
  wire[31:0] T117;
  wire[31:0] T118;
  wire T119;
  wire T120;
  wire T121;
  reg  wb_ctrl_wfd;
  wire T122;
  reg  mem_ctrl_wfd;
  wire T123;
  reg  ex_ctrl_wfd;
  wire T124;
  wire id_ctrl_wfd;
  wire T125;
  wire T126;
  wire[31:0] T127;
  wire T128;
  wire T129;
  wire[31:0] T130;
  wire T131;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire[31:0] T135;
  wire wb_dcache_miss;
  wire T136;
  reg  wb_ctrl_mem;
  wire T137;
  reg  mem_ctrl_mem;
  wire T138;
  reg  ex_ctrl_mem;
  wire T139;
  wire[31:0] T140;
  wire[31:0] T141;
  wire[31:0] T142;
  wire[31:0] T143;
  wire T144;
  wire[31:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[31:0] T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire[4:0] T155;
  wire[4:0] T156;
  wire[4:0] id_raddr3;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] id_raddr2;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire[4:0] T171;
  wire[4:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire id_ctrl_fp;
  wire T176;
  wire T177;
  wire[31:0] T178;
  wire T179;
  wire T180;
  wire[31:0] T181;
  wire T182;
  wire id_sboard_hazard;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[4:0] T187;
  wire[4:0] T188;
  wire T189;
  wire[31:0] T190;
  wire[31:0] T191;
  wire[31:0] T192;
  wire[31:0] T193;
  reg [31:0] R194;
  wire[31:0] T907;
  wire[31:0] T195;
  wire[31:0] T196;
  wire[31:0] T197;
  wire[31:0] T198;
  wire[31:0] T199;
  wire T200;
  wire wb_set_sboard;
  wire T201;
  reg  wb_ctrl_div;
  wire T202;
  reg  mem_ctrl_div;
  wire T203;
  reg  ex_ctrl_div;
  wire T204;
  wire id_ctrl_div;
  wire T205;
  wire[31:0] T206;
  wire T207;
  wire id_wen_not0;
  wire T208;
  wire id_ctrl_wxd;
  wire T209;
  wire T210;
  wire[31:0] T211;
  wire T212;
  wire T213;
  wire[31:0] T214;
  wire T215;
  wire T216;
  wire[31:0] T217;
  wire T218;
  wire T219;
  wire[31:0] T220;
  wire T221;
  wire T222;
  wire[31:0] T223;
  wire T224;
  wire T225;
  wire[31:0] T226;
  wire T227;
  wire T228;
  wire[31:0] T229;
  wire T230;
  wire[31:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[4:0] T237;
  wire[4:0] T238;
  wire T239;
  wire id_renx2_not0;
  wire T240;
  wire id_ctrl_rxs2;
  wire T241;
  wire T242;
  wire[31:0] T243;
  wire T244;
  wire T245;
  wire[31:0] T246;
  wire T247;
  wire T248;
  wire[31:0] T249;
  wire T250;
  wire[31:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[4:0] T256;
  wire[4:0] T257;
  wire T258;
  wire id_renx1_not0;
  wire T259;
  wire id_ctrl_rxs1;
  wire T260;
  wire T261;
  wire[31:0] T262;
  wire T263;
  wire T264;
  wire[31:0] T265;
  wire T266;
  wire T267;
  wire[31:0] T268;
  wire T269;
  wire T270;
  wire[31:0] T271;
  wire T272;
  wire T273;
  wire[31:0] T274;
  wire T275;
  wire T276;
  wire[31:0] T277;
  wire T278;
  wire[31:0] T279;
  wire T280;
  wire id_wb_hazard;
  wire T281;
  wire fp_data_hazard_wb;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire data_hazard_wb;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  reg  wb_ctrl_wxd;
  wire T302;
  reg  mem_ctrl_wxd;
  wire T303;
  reg  ex_ctrl_wxd;
  wire T304;
  wire T305;
  wire id_mem_hazard;
  wire T306;
  wire fp_data_hazard_mem;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire mem_cannot_bypass;
  wire T319;
  reg  mem_ctrl_fp;
  wire T320;
  reg  ex_ctrl_fp;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  reg  mem_mem_cmd_bh;
  wire T325;
  wire ex_slow_bypass;
  wire T326;
  wire T327;
  reg [3:0] ex_ctrl_mem_type;
  wire[3:0] T328;
  wire[3:0] id_ctrl_mem_type;
  wire[3:0] T329;
  wire[2:0] T330;
  wire[1:0] T331;
  wire T332;
  wire T333;
  wire[31:0] T334;
  wire T335;
  wire T336;
  wire[31:0] T337;
  wire T338;
  wire T339;
  wire[31:0] T340;
  wire T341;
  wire[31:0] T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  reg [4:0] ex_ctrl_mem_cmd;
  wire[4:0] T351;
  wire[4:0] id_ctrl_mem_cmd;
  wire[4:0] T352;
  wire[3:0] T353;
  wire[2:0] T354;
  wire[1:0] T355;
  wire T356;
  wire T357;
  wire[31:0] T358;
  wire T359;
  wire T360;
  wire[31:0] T361;
  wire T362;
  wire T363;
  wire[31:0] T364;
  wire T365;
  wire[31:0] T366;
  wire T367;
  wire T368;
  wire[31:0] T369;
  wire T370;
  wire[31:0] T371;
  wire T372;
  wire T373;
  wire[31:0] T374;
  wire T375;
  wire T376;
  wire[31:0] T377;
  wire T378;
  wire[31:0] T379;
  wire T380;
  reg [1:0] mem_ctrl_csr;
  wire[1:0] T381;
  reg [1:0] ex_ctrl_csr;
  wire[1:0] T382;
  wire data_hazard_mem;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  reg  mem_reg_valid;
  wire T391;
  wire ctrl_killx;
  wire T392;
  wire T393;
  reg  ex_reg_valid;
  wire T394;
  wire T395;
  wire replay_ex;
  wire T396;
  wire replay_ex_load_use;
  reg  ex_reg_load_use;
  wire T397;
  wire id_load_use;
  wire T398;
  wire T399;
  wire replay_ex_structural;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire take_pc;
  wire take_pc_mem;
  wire T404;
  reg  mem_reg_flush_pipe;
  wire T405;
  reg  ex_reg_flush_pipe;
  wire T406;
  wire T407;
  wire mem_misprediction;
  wire T408;
  reg  mem_ctrl_jal;
  wire T409;
  reg  ex_ctrl_jal;
  wire T410;
  wire id_ctrl_jal;
  wire T411;
  wire[31:0] T412;
  wire T413;
  reg  mem_ctrl_jalr;
  wire T414;
  reg  ex_ctrl_jalr;
  wire T415;
  wire id_ctrl_jalr;
  wire T416;
  wire[31:0] T417;
  reg  mem_ctrl_branch;
  wire T418;
  reg  ex_ctrl_branch;
  wire T419;
  wire id_ctrl_branch;
  wire T420;
  wire[31:0] T421;
  wire T422;
  wire id_ex_hazard;
  wire T423;
  wire fp_data_hazard_ex;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire ex_cannot_bypass;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire data_hazard_ex;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire ctrl_killm;
  wire T453;
  wire fpu_kill_mem;
  wire T454;
  wire T455;
  wire killm_common;
  wire T456;
  wire T457;
  reg  mem_reg_xcpt;
  wire T458;
  wire T459;
  wire T614;
  wire ex_xcpt;
  wire T460;
  wire T461;
  reg  ex_reg_xcpt;
  wire T462;
  wire T463;
  wire T610;
  wire id_xcpt;
  wire T464;
  wire T465;
  wire T466;
  wire id_ctrl_scall;
  wire T467;
  wire[31:0] T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire id_csr_fp;
  wire T473;
  wire[11:0] T474;
  wire T475;
  wire T476;
  wire T477;
  wire id_ctrl_sret;
  wire T478;
  wire[31:0] T479;
  wire T480;
  wire id_csr_privileged;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire[1:0] T486;
  wire T487;
  wire T488;
  wire[1:0] T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[1:0] T494;
  wire T495;
  wire T496;
  wire[1:0] T497;
  wire T498;
  wire T499;
  wire[1:0] T500;
  wire T501;
  wire T502;
  wire id_csr_invalid;
  wire T503;
  reg  T504;
  wire T506;
  wire id_ctrl_legal;
  wire T507;
  wire T508;
  wire[31:0] T509;
  wire T510;
  wire T511;
  wire[31:0] T512;
  wire T513;
  wire T514;
  wire[31:0] T515;
  wire T516;
  wire T517;
  wire[31:0] T518;
  wire T519;
  wire T520;
  wire[31:0] T521;
  wire T522;
  wire T523;
  wire[31:0] T524;
  wire T525;
  wire T526;
  wire[31:0] T527;
  wire T528;
  wire T529;
  wire[31:0] T530;
  wire T531;
  wire T532;
  wire[31:0] T533;
  wire T534;
  wire T535;
  wire[31:0] T536;
  wire T537;
  wire T538;
  wire[31:0] T539;
  wire T540;
  wire T541;
  wire[31:0] T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire[31:0] T547;
  wire T548;
  wire T549;
  wire[31:0] T550;
  wire T551;
  wire T552;
  wire[31:0] T553;
  wire T554;
  wire T555;
  wire[31:0] T556;
  wire T557;
  wire T558;
  wire[31:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[31:0] T563;
  wire T564;
  wire T565;
  wire T566;
  wire[31:0] T567;
  wire T568;
  wire T569;
  wire[31:0] T570;
  wire T571;
  wire T572;
  wire[31:0] T573;
  wire T574;
  wire T575;
  wire[31:0] T576;
  wire T577;
  wire T578;
  wire[31:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire[31:0] T583;
  wire T584;
  wire T585;
  wire[31:0] T586;
  wire T587;
  wire T588;
  wire[31:0] T589;
  wire T590;
  wire T591;
  wire[31:0] T592;
  wire T593;
  wire T594;
  wire[31:0] T595;
  wire T596;
  wire T597;
  wire[31:0] T598;
  wire T599;
  wire T600;
  wire[31:0] T601;
  wire T602;
  wire T603;
  wire[31:0] T604;
  wire T605;
  wire T606;
  wire[31:0] T607;
  wire T608;
  wire T609;
  reg  ex_reg_xcpt_interrupt;
  wire T611;
  wire T612;
  wire T613;
  wire T615;
  wire dcache_kill_mem;
  wire T616;
  reg  wb_reg_valid;
  wire T617;
  wire replay_wb_common;
  wire T618;
  reg  wb_reg_replay;
  wire T619;
  wire T620;
  wire replay_mem;
  wire T621;
  reg  mem_reg_replay;
  wire T622;
  wire T623;
  wire mem_xcpt;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  reg  mem_reg_xcpt_interrupt;
  wire T636;
  wire T637;
  wire wb_rocc_val;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  reg  wb_ctrl_fence_i;
  wire T645;
  reg  mem_ctrl_fence_i;
  wire T646;
  reg  ex_ctrl_fence_i;
  wire T647;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T648;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T649;
  wire T650;
  wire T651;
  reg  ex_reg_btb_hit;
  wire T652;
  reg [6:0] mem_reg_btb_resp_bht_history;
  wire[6:0] T653;
  reg [6:0] ex_reg_btb_resp_bht_history;
  wire[6:0] T654;
  reg [5:0] mem_reg_btb_resp_entry;
  wire[5:0] T655;
  reg [5:0] ex_reg_btb_resp_entry;
  wire[5:0] T656;
  reg [42:0] mem_reg_btb_resp_target;
  wire[42:0] T657;
  reg [42:0] ex_reg_btb_resp_target;
  wire[42:0] T658;
  reg  mem_reg_btb_resp_bridx;
  wire T659;
  reg  ex_reg_btb_resp_bridx;
  wire T660;
  reg  mem_reg_btb_resp_mask;
  wire T661;
  reg  ex_reg_btb_resp_mask;
  wire T662;
  reg  mem_reg_btb_resp_taken;
  wire T663;
  reg  ex_reg_btb_resp_taken;
  wire T664;
  reg  mem_reg_btb_hit;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  reg [63:0] wb_reg_cause;
  wire[63:0] T685;
  wire[63:0] mem_cause;
  wire[63:0] T908;
  wire[3:0] T686;
  wire[3:0] T687;
  wire[3:0] T688;
  reg [63:0] mem_reg_cause;
  wire[63:0] T689;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T690;
  wire[63:0] id_cause;
  wire[63:0] T909;
  wire[3:0] T691;
  wire[3:0] T692;
  wire[3:0] T693;
  wire[3:0] T694;
  wire[3:0] T695;
  wire[3:0] T696;
  wire[3:0] T697;
  wire[63:0] id_interrupt_cause;
  wire[63:0] T698;
  wire[63:0] T699;
  wire[63:0] T700;
  wire[63:0] T701;
  wire[63:0] T702;
  wire[63:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire[1:0] T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[1:0] T720;
  wire[1:0] T721;
  wire[1:0] T722;
  wire T723;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  reg  wb_ctrl_sret;
  wire T743;
  reg  mem_ctrl_sret;
  wire T744;
  reg  ex_ctrl_sret;
  wire T745;
  wire[2:0] T910;
  wire[1:0] T746;
  reg [1:0] wb_ctrl_csr;
  wire[1:0] T747;
  reg  mem_ctrl_amo;
  wire T748;
  reg  ex_ctrl_amo;
  wire T749;
  reg  mem_ctrl_fence;
  wire T750;
  reg  ex_ctrl_fence;
  wire T751;
  reg  mem_ctrl_scall;
  wire T752;
  reg  ex_ctrl_scall;
  wire T753;
  reg  mem_ctrl_rfs3;
  wire T754;
  reg  ex_ctrl_rfs3;
  wire T755;
  wire id_ctrl_rfs3;
  reg  mem_ctrl_rfs2;
  wire T756;
  reg  ex_ctrl_rfs2;
  wire T757;
  wire id_ctrl_rfs2;
  wire T758;
  wire T759;
  wire T760;
  wire[31:0] T761;
  wire T762;
  wire[31:0] T763;
  reg  mem_ctrl_rfs1;
  wire T764;
  reg  ex_ctrl_rfs1;
  wire T765;
  wire id_ctrl_rfs1;
  wire T766;
  wire T767;
  wire T768;
  wire[31:0] T769;
  reg [3:0] mem_ctrl_mem_type;
  wire[3:0] T770;
  reg [4:0] mem_ctrl_mem_cmd;
  wire[4:0] T771;
  reg [3:0] mem_ctrl_alu_fn;
  wire[3:0] T772;
  reg [3:0] ex_ctrl_alu_fn;
  wire[3:0] T773;
  wire[3:0] id_ctrl_alu_fn;
  wire[3:0] T774;
  wire[2:0] T775;
  wire[1:0] T776;
  wire T777;
  wire T778;
  wire[31:0] T779;
  wire T780;
  wire T781;
  wire[31:0] T782;
  wire T783;
  wire[31:0] T784;
  wire T785;
  wire T786;
  wire[31:0] T787;
  wire T788;
  wire T789;
  wire[31:0] T790;
  wire T791;
  wire T792;
  wire[31:0] T793;
  wire T794;
  wire T795;
  wire[31:0] T796;
  wire T797;
  wire[31:0] T798;
  wire T799;
  wire T800;
  wire[31:0] T801;
  wire T802;
  wire T803;
  wire[31:0] T804;
  wire T805;
  wire T806;
  wire[31:0] T807;
  wire T808;
  wire[31:0] T809;
  wire T810;
  wire T811;
  wire[31:0] T812;
  wire T813;
  wire T814;
  wire T815;
  wire[31:0] T816;
  wire T817;
  wire[31:0] T818;
  reg  mem_ctrl_alu_dw;
  wire T819;
  reg  ex_ctrl_alu_dw;
  wire T820;
  wire id_ctrl_alu_dw;
  wire T821;
  wire T822;
  wire[31:0] T823;
  wire T824;
  wire[31:0] T825;
  reg [2:0] mem_ctrl_sel_imm;
  wire[2:0] T826;
  reg [2:0] ex_ctrl_sel_imm;
  wire[2:0] T827;
  wire[2:0] id_ctrl_sel_imm;
  wire[2:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire[31:0] T832;
  wire T833;
  wire[31:0] T834;
  wire T835;
  wire T836;
  wire[31:0] T837;
  wire T838;
  wire T839;
  wire[31:0] T840;
  wire T841;
  wire T842;
  wire[31:0] T843;
  wire T844;
  wire T845;
  wire[31:0] T846;
  wire T847;
  wire[31:0] T848;
  reg [1:0] mem_ctrl_sel_alu1;
  wire[1:0] T849;
  reg [1:0] ex_ctrl_sel_alu1;
  wire[1:0] T850;
  wire[1:0] id_ctrl_sel_alu1;
  wire[1:0] T851;
  wire T852;
  wire T853;
  wire[31:0] T854;
  wire T855;
  wire T856;
  wire[31:0] T857;
  wire T858;
  wire T859;
  wire T860;
  wire[31:0] T861;
  wire T862;
  wire[31:0] T863;
  wire T864;
  wire T865;
  wire[31:0] T866;
  wire T867;
  wire[31:0] T868;
  reg [1:0] mem_ctrl_sel_alu2;
  wire[1:0] T869;
  reg [1:0] ex_ctrl_sel_alu2;
  wire[1:0] T870;
  wire[1:0] id_ctrl_sel_alu2;
  wire[1:0] T871;
  wire T872;
  wire T873;
  wire[31:0] T874;
  wire T875;
  wire T876;
  wire T877;
  wire[31:0] T878;
  wire T879;
  wire T880;
  wire[31:0] T881;
  wire T882;
  wire[31:0] T883;
  wire T884;
  wire T885;
  wire[31:0] T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire[31:0] T891;
  reg  mem_ctrl_rxs1;
  wire T892;
  reg  ex_ctrl_rxs1;
  wire T893;
  reg  mem_ctrl_rxs2;
  wire T894;
  reg  ex_ctrl_rxs2;
  wire T895;
  reg  mem_ctrl_legal;
  wire T896;
  reg  ex_ctrl_legal;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire[2:0] T911;
  wire[1:0] T901;
  wire[1:0] T902;
  wire[1:0] T903;
  wire T904;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wb_reg_xcpt = {1{$random}};
    wb_ctrl_rocc = {1{$random}};
    mem_ctrl_rocc = {1{$random}};
    ex_ctrl_rocc = {1{$random}};
    id_reg_fence = {1{$random}};
    R112 = {1{$random}};
    wb_ctrl_wfd = {1{$random}};
    mem_ctrl_wfd = {1{$random}};
    ex_ctrl_wfd = {1{$random}};
    wb_ctrl_mem = {1{$random}};
    mem_ctrl_mem = {1{$random}};
    ex_ctrl_mem = {1{$random}};
    R194 = {1{$random}};
    wb_ctrl_div = {1{$random}};
    mem_ctrl_div = {1{$random}};
    ex_ctrl_div = {1{$random}};
    wb_ctrl_wxd = {1{$random}};
    mem_ctrl_wxd = {1{$random}};
    ex_ctrl_wxd = {1{$random}};
    mem_ctrl_fp = {1{$random}};
    ex_ctrl_fp = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_ctrl_mem_type = {1{$random}};
    ex_ctrl_mem_cmd = {1{$random}};
    mem_ctrl_csr = {1{$random}};
    ex_ctrl_csr = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_reg_flush_pipe = {1{$random}};
    ex_reg_flush_pipe = {1{$random}};
    mem_ctrl_jal = {1{$random}};
    ex_ctrl_jal = {1{$random}};
    mem_ctrl_jalr = {1{$random}};
    ex_ctrl_jalr = {1{$random}};
    mem_ctrl_branch = {1{$random}};
    ex_ctrl_branch = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    wb_reg_valid = {1{$random}};
    wb_reg_replay = {1{$random}};
    mem_reg_replay = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    wb_ctrl_fence_i = {1{$random}};
    mem_ctrl_fence_i = {1{$random}};
    ex_ctrl_fence_i = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_bridx = {1{$random}};
    ex_reg_btb_resp_bridx = {1{$random}};
    mem_reg_btb_resp_mask = {1{$random}};
    ex_reg_btb_resp_mask = {1{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_ctrl_sret = {1{$random}};
    mem_ctrl_sret = {1{$random}};
    ex_ctrl_sret = {1{$random}};
    wb_ctrl_csr = {1{$random}};
    mem_ctrl_amo = {1{$random}};
    ex_ctrl_amo = {1{$random}};
    mem_ctrl_fence = {1{$random}};
    ex_ctrl_fence = {1{$random}};
    mem_ctrl_scall = {1{$random}};
    ex_ctrl_scall = {1{$random}};
    mem_ctrl_rfs3 = {1{$random}};
    ex_ctrl_rfs3 = {1{$random}};
    mem_ctrl_rfs2 = {1{$random}};
    ex_ctrl_rfs2 = {1{$random}};
    mem_ctrl_rfs1 = {1{$random}};
    ex_ctrl_rfs1 = {1{$random}};
    mem_ctrl_mem_type = {1{$random}};
    mem_ctrl_mem_cmd = {1{$random}};
    mem_ctrl_alu_fn = {1{$random}};
    ex_ctrl_alu_fn = {1{$random}};
    mem_ctrl_alu_dw = {1{$random}};
    ex_ctrl_alu_dw = {1{$random}};
    mem_ctrl_sel_imm = {1{$random}};
    ex_ctrl_sel_imm = {1{$random}};
    mem_ctrl_sel_alu1 = {1{$random}};
    ex_ctrl_sel_alu1 = {1{$random}};
    mem_ctrl_sel_alu2 = {1{$random}};
    ex_ctrl_sel_alu2 = {1{$random}};
    mem_ctrl_rxs1 = {1{$random}};
    ex_ctrl_rxs1 = {1{$random}};
    mem_ctrl_rxs2 = {1{$random}};
    ex_ctrl_rxs2 = {1{$random}};
    mem_ctrl_legal = {1{$random}};
    ex_ctrl_legal = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rocc_exception = T0;
  assign T0 = wb_reg_xcpt & io_dpath_status_er;
  assign T1 = mem_xcpt & T2;
  assign T2 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T3;
  assign T3 = T4 | io_dpath_sret;
  assign T4 = replay_wb | wb_reg_xcpt;
  assign replay_wb = replay_wb_common | T5;
  assign T5 = T7 & T6;
  assign T6 = io_rocc_cmd_ready ^ 1'h1;
  assign T7 = wb_reg_valid & wb_ctrl_rocc;
  assign T8 = T452 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign T9 = T451 ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign T10 = T11 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign id_ctrl_rocc = 1'h0;
  assign T11 = ctrl_killd ^ 1'h1;
  assign ctrl_killd = T12;
  assign T12 = T43 | ctrl_draind;
  assign ctrl_draind = io_dpath_status_ei & id_interrupt_unmasked;
  assign id_interrupt_unmasked = T16 | T13;
  assign T13 = T15 & T14;
  assign T14 = io_dpath_status_ip[3'h7:3'h7];
  assign T15 = io_dpath_status_im[3'h7:3'h7];
  assign T16 = T20 | T17;
  assign T17 = T19 & T18;
  assign T18 = io_dpath_status_ip[3'h6:3'h6];
  assign T19 = io_dpath_status_im[3'h6:3'h6];
  assign T20 = T24 | T21;
  assign T21 = T23 & T22;
  assign T22 = io_dpath_status_ip[3'h5:3'h5];
  assign T23 = io_dpath_status_im[3'h5:3'h5];
  assign T24 = T28 | T25;
  assign T25 = T27 & T26;
  assign T26 = io_dpath_status_ip[3'h4:3'h4];
  assign T27 = io_dpath_status_im[3'h4:3'h4];
  assign T28 = T32 | T29;
  assign T29 = T31 & T30;
  assign T30 = io_dpath_status_ip[2'h3:2'h3];
  assign T31 = io_dpath_status_im[2'h3:2'h3];
  assign T32 = T36 | T33;
  assign T33 = T35 & T34;
  assign T34 = io_dpath_status_ip[2'h2:2'h2];
  assign T35 = io_dpath_status_im[2'h2:2'h2];
  assign T36 = T40 | T37;
  assign T37 = T39 & T38;
  assign T38 = io_dpath_status_ip[1'h1:1'h1];
  assign T39 = io_dpath_status_im[1'h1:1'h1];
  assign T40 = T42 & T41;
  assign T41 = io_dpath_status_ip[1'h0:1'h0];
  assign T42 = io_dpath_status_im[1'h0:1'h0];
  assign T43 = T449 | ctrl_stalld;
  assign ctrl_stalld = T100 | id_do_fence;
  assign id_do_fence = id_mem_busy & T44;
  assign T44 = T62 | id_csr_flush;
  assign id_csr_flush = T51 & T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T49 | T47;
  assign T47 = T48 == 12'h400;
  assign T48 = id_csr_addr & 12'hc2d;
  assign id_csr_addr = io_dpath_inst[5'h1f:5'h14];
  assign T49 = T50 == 12'h400;
  assign T50 = id_csr_addr & 12'hc2e;
  assign T51 = id_csr_en & id_csr_wen;
  assign id_csr_wen = T61 | T52;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T60 | T54;
  assign T54 = 2'h3 == id_ctrl_csr;
  assign id_ctrl_csr = T55;
  assign T55 = {T58, T56};
  assign T56 = T57 == 32'h1070;
  assign T57 = io_dpath_inst & 32'h1070;
  assign T58 = T59 == 32'h2070;
  assign T59 = io_dpath_inst & 32'h2070;
  assign T60 = 2'h2 == id_ctrl_csr;
  assign T61 = id_raddr1 != 5'h0;
  assign id_raddr1 = io_dpath_inst[5'h13:4'hf];
  assign id_csr_en = id_ctrl_csr != 2'h0;
  assign T62 = T95 | T63;
  assign T63 = id_reg_fence & T64;
  assign T64 = id_ctrl_mem | id_ctrl_rocc;
  assign id_ctrl_mem = T65;
  assign T65 = T68 | T66;
  assign T66 = T67 == 32'h1000202f;
  assign T67 = io_dpath_inst & 32'hf9f0607f;
  assign T68 = T71 | T69;
  assign T69 = T70 == 32'h800202f;
  assign T70 = io_dpath_inst & 32'he800607f;
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h202f;
  assign T73 = io_dpath_inst & 32'h1800607f;
  assign T74 = T77 | T75;
  assign T75 = T76 == 32'h2003;
  assign T76 = io_dpath_inst & 32'h605b;
  assign T77 = T80 | T78;
  assign T78 = T79 == 32'h57;
  assign T79 = io_dpath_inst & 32'h607f;
  assign T80 = T83 | T81;
  assign T81 = T82 == 32'h3;
  assign T82 = io_dpath_inst & 32'h107f;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h3;
  assign T85 = io_dpath_inst & 32'h207f;
  assign T86 = T87 == 32'h3;
  assign T87 = io_dpath_inst & 32'h405f;
  assign T905 = reset ? 1'h0 : T88;
  assign T88 = id_fence_next | T89;
  assign T89 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_ctrl_fence | T90;
  assign T90 = id_ctrl_amo & id_amo_rl;
  assign id_amo_rl = io_dpath_inst[5'h19:5'h19];
  assign id_ctrl_amo = T91;
  assign T91 = T92 == 32'h2008;
  assign T92 = io_dpath_inst & 32'h6048;
  assign id_ctrl_fence = T93;
  assign T93 = T94 == 32'h8;
  assign T94 = io_dpath_inst & 32'h3058;
  assign T95 = T98 | id_ctrl_fence_i;
  assign id_ctrl_fence_i = T96;
  assign T96 = T97 == 32'h1008;
  assign T97 = io_dpath_inst & 32'h3058;
  assign T98 = id_ctrl_amo & id_amo_aq;
  assign id_amo_aq = io_dpath_inst[5'h1a:5'h1a];
  assign id_mem_busy = T99 | io_dmem_req_valid;
  assign T99 = io_dmem_ordered ^ 1'h1;
  assign T100 = T103 | T101;
  assign T101 = id_ctrl_mem & T102;
  assign T102 = io_dmem_req_ready ^ 1'h1;
  assign T103 = T182 | T104;
  assign T104 = id_ctrl_fp & id_stall_fpu;
  assign id_stall_fpu = T150 | T105;
  assign T105 = io_fpu_dec_wen & T106;
  assign T106 = T111 & T107;
  assign T107 = T108 - 1'h1;
  assign T108 = 1'h1 << T109;
  assign T109 = T110 + 5'h1;
  assign T110 = id_waddr - id_waddr;
  assign id_waddr = io_dpath_inst[4'hb:3'h7];
  assign T111 = R112 >> id_waddr;
  assign T906 = reset ? 32'h0 : T113;
  assign T113 = T149 ? T145 : T114;
  assign T114 = T144 ? T140 : T115;
  assign T115 = T119 ? T116 : R112;
  assign T116 = R112 | T117;
  assign T117 = T119 ? T118 : 32'h0;
  assign T118 = 1'h1 << io_dpath_wb_waddr;
  assign T119 = T120 & io_dpath_retire;
  assign T120 = T121 | io_fpu_sboard_set;
  assign T121 = wb_dcache_miss & wb_ctrl_wfd;
  assign T122 = T452 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign T123 = T451 ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign T124 = T11 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign id_ctrl_wfd = T125;
  assign T125 = T128 | T126;
  assign T126 = T127 == 32'h10000040;
  assign T127 = io_dpath_inst & 32'h10000064;
  assign T128 = T131 | T129;
  assign T129 = T130 == 32'h40;
  assign T130 = io_dpath_inst & 32'h70;
  assign T131 = T134 | T132;
  assign T132 = T133 == 32'h40;
  assign T133 = io_dpath_inst & 32'h80000064;
  assign T134 = T135 == 32'h4;
  assign T135 = io_dpath_inst & 32'h3c;
  assign wb_dcache_miss = wb_ctrl_mem & T136;
  assign T136 = io_dmem_resp_valid ^ 1'h1;
  assign T137 = T452 ? mem_ctrl_mem : wb_ctrl_mem;
  assign T138 = T451 ? ex_ctrl_mem : mem_ctrl_mem;
  assign T139 = T11 ? id_ctrl_mem : ex_ctrl_mem;
  assign T140 = T116 & T141;
  assign T141 = ~ T142;
  assign T142 = io_dpath_fp_sboard_clr ? T143 : 32'h0;
  assign T143 = 1'h1 << io_dpath_fp_sboard_clra;
  assign T144 = T119 | io_dpath_fp_sboard_clr;
  assign T145 = T140 & T146;
  assign T146 = ~ T147;
  assign T147 = io_fpu_sboard_clr ? T148 : 32'h0;
  assign T148 = 1'h1 << io_fpu_sboard_clra;
  assign T149 = T144 | io_fpu_sboard_clr;
  assign T150 = T158 | T151;
  assign T151 = io_fpu_dec_ren3 & T152;
  assign T152 = T157 & T153;
  assign T153 = T154 - 1'h1;
  assign T154 = 1'h1 << T155;
  assign T155 = T156 + 5'h1;
  assign T156 = id_raddr3 - id_raddr3;
  assign id_raddr3 = io_dpath_inst[5'h1f:5'h1b];
  assign T157 = R112 >> id_raddr3;
  assign T158 = T166 | T159;
  assign T159 = io_fpu_dec_ren2 & T160;
  assign T160 = T165 & T161;
  assign T161 = T162 - 1'h1;
  assign T162 = 1'h1 << T163;
  assign T163 = T164 + 5'h1;
  assign T164 = id_raddr2 - id_raddr2;
  assign id_raddr2 = io_dpath_inst[5'h18:5'h14];
  assign T165 = R112 >> id_raddr2;
  assign T166 = T174 | T167;
  assign T167 = io_fpu_dec_ren1 & T168;
  assign T168 = T173 & T169;
  assign T169 = T170 - 1'h1;
  assign T170 = 1'h1 << T171;
  assign T171 = T172 + 5'h1;
  assign T172 = id_raddr1 - id_raddr1;
  assign T173 = R112 >> id_raddr1;
  assign T174 = id_csr_en & T175;
  assign T175 = io_fpu_fcsr_rdy ^ 1'h1;
  assign id_ctrl_fp = T176;
  assign T176 = T179 | T177;
  assign T177 = T178 == 32'h40;
  assign T178 = io_dpath_inst & 32'h64;
  assign T179 = T180 | T129;
  assign T180 = T181 == 32'h4;
  assign T181 = io_dpath_inst & 32'h5c;
  assign T182 = T280 | id_sboard_hazard;
  assign id_sboard_hazard = T232 | T183;
  assign T183 = id_wen_not0 & T184;
  assign T184 = T189 & T185;
  assign T185 = T186 - 1'h1;
  assign T186 = 1'h1 << T187;
  assign T187 = T188 + 5'h1;
  assign T188 = id_waddr - id_waddr;
  assign T189 = T190 >> id_waddr;
  assign T190 = R194 & T191;
  assign T191 = ~ T192;
  assign T192 = io_dpath_ll_wen ? T193 : 32'h0;
  assign T193 = 1'h1 << io_dpath_ll_waddr;
  assign T907 = reset ? 32'h0 : T195;
  assign T195 = T207 ? T197 : T196;
  assign T196 = io_dpath_ll_wen ? T190 : R194;
  assign T197 = T190 | T198;
  assign T198 = T200 ? T199 : 32'h0;
  assign T199 = 1'h1 << io_dpath_wb_waddr;
  assign T200 = wb_set_sboard & io_dpath_wb_wen;
  assign wb_set_sboard = T201 | wb_ctrl_rocc;
  assign T201 = wb_ctrl_div | wb_dcache_miss;
  assign T202 = T452 ? mem_ctrl_div : wb_ctrl_div;
  assign T203 = T451 ? ex_ctrl_div : mem_ctrl_div;
  assign T204 = T11 ? id_ctrl_div : ex_ctrl_div;
  assign id_ctrl_div = T205;
  assign T205 = T206 == 32'h2000030;
  assign T206 = io_dpath_inst & 32'h2000074;
  assign T207 = io_dpath_ll_wen | T200;
  assign id_wen_not0 = id_ctrl_wxd & T208;
  assign T208 = id_waddr != 5'h0;
  assign id_ctrl_wxd = T209;
  assign T209 = T212 | T210;
  assign T210 = T211 == 32'h80000010;
  assign T211 = io_dpath_inst & 32'h90000034;
  assign T212 = T215 | T213;
  assign T213 = T214 == 32'h2030;
  assign T214 = io_dpath_inst & 32'h2030;
  assign T215 = T218 | T216;
  assign T216 = T217 == 32'h1030;
  assign T217 = io_dpath_inst & 32'h1030;
  assign T218 = T221 | T219;
  assign T219 = T220 == 32'h28;
  assign T220 = io_dpath_inst & 32'h28;
  assign T221 = T224 | T222;
  assign T222 = T223 == 32'h24;
  assign T223 = io_dpath_inst & 32'h2024;
  assign T224 = T227 | T225;
  assign T225 = T226 == 32'h14;
  assign T226 = io_dpath_inst & 32'h1014;
  assign T227 = T230 | T228;
  assign T228 = T229 == 32'h10;
  assign T229 = io_dpath_inst & 32'h50;
  assign T230 = T231 == 32'h0;
  assign T231 = io_dpath_inst & 32'h64;
  assign T232 = T252 | T233;
  assign T233 = id_renx2_not0 & T234;
  assign T234 = T239 & T235;
  assign T235 = T236 - 1'h1;
  assign T236 = 1'h1 << T237;
  assign T237 = T238 + 5'h1;
  assign T238 = id_raddr2 - id_raddr2;
  assign T239 = T190 >> id_raddr2;
  assign id_renx2_not0 = id_ctrl_rxs2 & T240;
  assign T240 = id_raddr2 != 5'h0;
  assign id_ctrl_rxs2 = T241;
  assign T241 = T244 | T242;
  assign T242 = T243 == 32'h2008;
  assign T243 = io_dpath_inst & 32'h2048;
  assign T244 = T247 | T245;
  assign T245 = T246 == 32'h1054;
  assign T246 = io_dpath_inst & 32'h1054;
  assign T247 = T250 | T248;
  assign T248 = T249 == 32'h20;
  assign T249 = io_dpath_inst & 32'h34;
  assign T250 = T251 == 32'h20;
  assign T251 = io_dpath_inst & 32'h64;
  assign T252 = id_renx1_not0 & T253;
  assign T253 = T258 & T254;
  assign T254 = T255 - 1'h1;
  assign T255 = 1'h1 << T256;
  assign T256 = T257 + 5'h1;
  assign T257 = id_raddr1 - id_raddr1;
  assign T258 = T190 >> id_raddr1;
  assign id_renx1_not0 = id_ctrl_rxs1 & T259;
  assign T259 = id_raddr1 != 5'h0;
  assign id_ctrl_rxs1 = T260;
  assign T260 = T263 | T261;
  assign T261 = T262 == 32'h90000010;
  assign T262 = io_dpath_inst & 32'h90000034;
  assign T263 = T266 | T264;
  assign T264 = T265 == 32'h2020;
  assign T265 = io_dpath_inst & 32'h6024;
  assign T266 = T269 | T267;
  assign T267 = T268 == 32'h2000;
  assign T268 = io_dpath_inst & 32'h2050;
  assign T269 = T272 | T270;
  assign T270 = T271 == 32'h1020;
  assign T271 = io_dpath_inst & 32'h5024;
  assign T272 = T275 | T273;
  assign T273 = T274 == 32'h54;
  assign T274 = io_dpath_inst & 32'h54;
  assign T275 = T278 | T276;
  assign T276 = T277 == 32'h20;
  assign T277 = io_dpath_inst & 32'h38;
  assign T278 = T279 == 32'h0;
  assign T279 = io_dpath_inst & 32'h44;
  assign T280 = T305 | id_wb_hazard;
  assign id_wb_hazard = wb_reg_valid & T281;
  assign T281 = T293 | fp_data_hazard_wb;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T282;
  assign T282 = T285 | T283;
  assign T283 = io_fpu_dec_wen & T284;
  assign T284 = id_waddr == io_dpath_wb_waddr;
  assign T285 = T288 | T286;
  assign T286 = io_fpu_dec_ren3 & T287;
  assign T287 = id_raddr3 == io_dpath_wb_waddr;
  assign T288 = T291 | T289;
  assign T289 = io_fpu_dec_ren2 & T290;
  assign T290 = id_raddr2 == io_dpath_wb_waddr;
  assign T291 = io_fpu_dec_ren1 & T292;
  assign T292 = id_raddr1 == io_dpath_wb_waddr;
  assign T293 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_ctrl_wxd & T294;
  assign T294 = T297 | T295;
  assign T295 = id_wen_not0 & T296;
  assign T296 = id_waddr == io_dpath_wb_waddr;
  assign T297 = T300 | T298;
  assign T298 = id_renx2_not0 & T299;
  assign T299 = id_raddr2 == io_dpath_wb_waddr;
  assign T300 = id_renx1_not0 & T301;
  assign T301 = id_raddr1 == io_dpath_wb_waddr;
  assign T302 = T452 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign T303 = T451 ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign T304 = T11 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign T305 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = mem_reg_valid & T306;
  assign T306 = T318 | fp_data_hazard_mem;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T307;
  assign T307 = T310 | T308;
  assign T308 = io_fpu_dec_wen & T309;
  assign T309 = id_waddr == io_dpath_mem_waddr;
  assign T310 = T313 | T311;
  assign T311 = io_fpu_dec_ren3 & T312;
  assign T312 = id_raddr3 == io_dpath_mem_waddr;
  assign T313 = T316 | T314;
  assign T314 = io_fpu_dec_ren2 & T315;
  assign T315 = id_raddr2 == io_dpath_mem_waddr;
  assign T316 = io_fpu_dec_ren1 & T317;
  assign T317 = id_raddr1 == io_dpath_mem_waddr;
  assign T318 = data_hazard_mem & mem_cannot_bypass;
  assign mem_cannot_bypass = T319 | mem_ctrl_rocc;
  assign T319 = T322 | mem_ctrl_fp;
  assign T320 = T451 ? ex_ctrl_fp : mem_ctrl_fp;
  assign T321 = T11 ? id_ctrl_fp : ex_ctrl_fp;
  assign T322 = T323 | mem_ctrl_div;
  assign T323 = T380 | T324;
  assign T324 = mem_ctrl_mem & mem_mem_cmd_bh;
  assign T325 = T451 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T350 | T326;
  assign T326 = T343 | T327;
  assign T327 = 4'hf == ex_ctrl_mem_type;
  assign T328 = T11 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign id_ctrl_mem_type = T329;
  assign T329 = {T341, T330};
  assign T330 = {T338, T331};
  assign T331 = {T335, T332};
  assign T332 = T341 | T333;
  assign T333 = T334 == 32'h1000;
  assign T334 = io_dpath_inst & 32'h1000;
  assign T335 = T341 | T336;
  assign T336 = T337 == 32'h2000;
  assign T337 = io_dpath_inst & 32'h2000;
  assign T338 = T341 | T339;
  assign T339 = T340 == 32'h4000;
  assign T340 = io_dpath_inst & 32'h4000;
  assign T341 = T342 == 32'h40;
  assign T342 = io_dpath_inst & 32'h40;
  assign T343 = T345 | T344;
  assign T344 = 4'h5 == ex_ctrl_mem_type;
  assign T345 = T347 | T346;
  assign T346 = 4'h1 == ex_ctrl_mem_type;
  assign T347 = T349 | T348;
  assign T348 = 4'h4 == ex_ctrl_mem_type;
  assign T349 = 4'h0 == ex_ctrl_mem_type;
  assign T350 = ex_ctrl_mem_cmd == 5'h7;
  assign T351 = T11 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign id_ctrl_mem_cmd = T352;
  assign T352 = {1'h0, T353};
  assign T353 = {T378, T354};
  assign T354 = {T372, T355};
  assign T355 = {T367, T356};
  assign T356 = T359 | T357;
  assign T357 = T358 == 32'h20000020;
  assign T358 = io_dpath_inst & 32'h20000020;
  assign T359 = T362 | T360;
  assign T360 = T361 == 32'h18000020;
  assign T361 = io_dpath_inst & 32'h18000020;
  assign T362 = T365 | T363;
  assign T363 = T364 == 32'h1040;
  assign T364 = io_dpath_inst & 32'h1040;
  assign T365 = T366 == 32'h20;
  assign T366 = io_dpath_inst & 32'h28;
  assign T367 = T370 | T368;
  assign T368 = T369 == 32'h40000008;
  assign T369 = io_dpath_inst & 32'h40000008;
  assign T370 = T371 == 32'h10000008;
  assign T371 = io_dpath_inst & 32'h10000008;
  assign T372 = T375 | T373;
  assign T373 = T374 == 32'h80000008;
  assign T374 = io_dpath_inst & 32'h80000008;
  assign T375 = T376 | T370;
  assign T376 = T377 == 32'h8000008;
  assign T377 = io_dpath_inst & 32'h8000008;
  assign T378 = T379 == 32'h8;
  assign T379 = io_dpath_inst & 32'h18000008;
  assign T380 = mem_ctrl_csr != 2'h0;
  assign T381 = T451 ? ex_ctrl_csr : mem_ctrl_csr;
  assign T382 = T11 ? id_ctrl_csr : ex_ctrl_csr;
  assign data_hazard_mem = mem_ctrl_wxd & T383;
  assign T383 = T386 | T384;
  assign T384 = id_wen_not0 & T385;
  assign T385 = id_waddr == io_dpath_mem_waddr;
  assign T386 = T389 | T387;
  assign T387 = id_renx2_not0 & T388;
  assign T388 = id_raddr2 == io_dpath_mem_waddr;
  assign T389 = id_renx1_not0 & T390;
  assign T390 = id_raddr1 == io_dpath_mem_waddr;
  assign T391 = ctrl_killx ^ 1'h1;
  assign ctrl_killx = T392;
  assign T392 = T395 | T393;
  assign T393 = ex_reg_valid ^ 1'h1;
  assign T394 = ctrl_killd ^ 1'h1;
  assign T395 = take_pc | replay_ex;
  assign replay_ex = ex_reg_valid & T396;
  assign T396 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T397 = T11 ? id_load_use : ex_reg_load_use;
  assign id_load_use = T398;
  assign T398 = T399 & mem_ctrl_mem;
  assign T399 = mem_reg_valid & data_hazard_mem;
  assign replay_ex_structural = T402 | T400;
  assign T400 = ex_ctrl_div & T401;
  assign T401 = io_dpath_div_mul_rdy ^ 1'h1;
  assign T402 = ex_ctrl_mem & T403;
  assign T403 = io_dmem_req_ready ^ 1'h1;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = mem_reg_valid & T404;
  assign T404 = mem_misprediction | mem_reg_flush_pipe;
  assign T405 = T451 ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign T406 = T11 ? T407 : ex_reg_flush_pipe;
  assign T407 = id_ctrl_fence_i | id_csr_flush;
  assign mem_misprediction = T422 & T408;
  assign T408 = T413 | mem_ctrl_jal;
  assign T409 = T451 ? ex_ctrl_jal : mem_ctrl_jal;
  assign T410 = T11 ? id_ctrl_jal : ex_ctrl_jal;
  assign id_ctrl_jal = T411;
  assign T411 = T412 == 32'h68;
  assign T412 = io_dpath_inst & 32'h68;
  assign T413 = mem_ctrl_branch | mem_ctrl_jalr;
  assign T414 = T451 ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign T415 = T11 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign id_ctrl_jalr = T416;
  assign T416 = T417 == 32'h24;
  assign T417 = io_dpath_inst & 32'h203c;
  assign T418 = T451 ? ex_ctrl_branch : mem_ctrl_branch;
  assign T419 = T11 ? id_ctrl_branch : ex_ctrl_branch;
  assign id_ctrl_branch = T420;
  assign T420 = T421 == 32'h60;
  assign T421 = io_dpath_inst & 32'h74;
  assign T422 = io_dpath_mem_misprediction & mem_reg_valid;
  assign id_ex_hazard = ex_reg_valid & T423;
  assign T423 = T435 | fp_data_hazard_ex;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T424;
  assign T424 = T427 | T425;
  assign T425 = io_fpu_dec_wen & T426;
  assign T426 = id_waddr == io_dpath_ex_waddr;
  assign T427 = T430 | T428;
  assign T428 = io_fpu_dec_ren3 & T429;
  assign T429 = id_raddr3 == io_dpath_ex_waddr;
  assign T430 = T433 | T431;
  assign T431 = io_fpu_dec_ren2 & T432;
  assign T432 = id_raddr2 == io_dpath_ex_waddr;
  assign T433 = io_fpu_dec_ren1 & T434;
  assign T434 = id_raddr1 == io_dpath_ex_waddr;
  assign T435 = data_hazard_ex & ex_cannot_bypass;
  assign ex_cannot_bypass = T436 | ex_ctrl_rocc;
  assign T436 = T437 | ex_ctrl_fp;
  assign T437 = T438 | ex_ctrl_div;
  assign T438 = T439 | ex_ctrl_mem;
  assign T439 = T440 | ex_ctrl_jalr;
  assign T440 = ex_ctrl_csr != 2'h0;
  assign data_hazard_ex = ex_ctrl_wxd & T441;
  assign T441 = T444 | T442;
  assign T442 = id_wen_not0 & T443;
  assign T443 = id_waddr == io_dpath_ex_waddr;
  assign T444 = T447 | T445;
  assign T445 = id_renx2_not0 & T446;
  assign T446 = id_raddr2 == io_dpath_ex_waddr;
  assign T447 = id_renx1_not0 & T448;
  assign T448 = id_raddr1 == io_dpath_ex_waddr;
  assign T449 = T450 | take_pc;
  assign T450 = io_imem_resp_valid ^ 1'h1;
  assign T451 = ctrl_killx ^ 1'h1;
  assign T452 = ctrl_killm ^ 1'h1;
  assign ctrl_killm = T453;
  assign T453 = T455 | fpu_kill_mem;
  assign fpu_kill_mem = T454 & io_fpu_nack_mem;
  assign T454 = mem_reg_valid & mem_ctrl_fp;
  assign T455 = killm_common | mem_xcpt;
  assign killm_common = T457 | T456;
  assign T456 = mem_reg_valid ^ 1'h1;
  assign T457 = T615 | mem_reg_xcpt;
  assign T458 = T451 ? ex_xcpt : T459;
  assign T459 = T614 & ex_xcpt;
  assign T614 = ctrl_killx ^ 1'h1;
  assign ex_xcpt = T461 | T460;
  assign T460 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign T461 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T462 = T11 ? id_xcpt : T463;
  assign T463 = T610 & id_xcpt;
  assign T610 = ctrl_killd ^ 1'h1;
  assign id_xcpt = T466 | T464;
  assign T464 = id_ctrl_rocc & T465;
  assign T465 = io_dpath_status_er ^ 1'h1;
  assign T466 = T469 | id_ctrl_scall;
  assign id_ctrl_scall = T467;
  assign T467 = T468 == 32'h70;
  assign T468 = io_dpath_inst & 32'h80003070;
  assign T469 = T475 | T470;
  assign T470 = T472 & T471;
  assign T471 = io_dpath_status_ef ^ 1'h1;
  assign T472 = id_ctrl_fp | id_csr_fp;
  assign id_csr_fp = id_csr_en & T473;
  assign T473 = T474 == 12'h0;
  assign T474 = id_csr_addr & 12'h480;
  assign T475 = T480 | T476;
  assign T476 = id_ctrl_sret & T477;
  assign T477 = io_dpath_status_s ^ 1'h1;
  assign id_ctrl_sret = T478;
  assign T478 = T479 == 32'h80000050;
  assign T479 = io_dpath_inst & 32'he0003054;
  assign T480 = T501 | id_csr_privileged;
  assign id_csr_privileged = id_csr_en & T481;
  assign T481 = T487 | T482;
  assign T482 = T483 & id_csr_wen;
  assign T483 = T485 & T484;
  assign T484 = io_dpath_status_s ^ 1'h1;
  assign T485 = T486 == 2'h1;
  assign T486 = id_csr_addr[4'h9:4'h8];
  assign T487 = T490 | T488;
  assign T488 = 2'h2 <= T489;
  assign T489 = id_csr_addr[4'h9:4'h8];
  assign T490 = T495 | T491;
  assign T491 = T493 & T492;
  assign T492 = io_dpath_status_s ^ 1'h1;
  assign T493 = T494 == 2'h1;
  assign T494 = id_csr_addr[4'hb:4'ha];
  assign T495 = T498 | T496;
  assign T496 = T497 == 2'h2;
  assign T497 = id_csr_addr[4'hb:4'ha];
  assign T498 = T499 & id_csr_wen;
  assign T499 = T500 == 2'h3;
  assign T500 = id_csr_addr[4'hb:4'ha];
  assign T501 = T608 | T502;
  assign T502 = T506 | id_csr_invalid;
  assign id_csr_invalid = id_csr_en & T503;
  assign T503 = T504 ^ 1'h1;
  always @(*) case (id_csr_addr)
    0: T504 = 1'h0;
    1: T504 = 1'h1;
    2: T504 = 1'h1;
    3: T504 = 1'h1;
    4: T504 = 1'h0;
    5: T504 = 1'h0;
    6: T504 = 1'h0;
    7: T504 = 1'h0;
    8: T504 = 1'h0;
    9: T504 = 1'h0;
    10: T504 = 1'h0;
    11: T504 = 1'h0;
    12: T504 = 1'h0;
    13: T504 = 1'h0;
    14: T504 = 1'h0;
    15: T504 = 1'h0;
    16: T504 = 1'h0;
    17: T504 = 1'h0;
    18: T504 = 1'h0;
    19: T504 = 1'h0;
    20: T504 = 1'h0;
    21: T504 = 1'h0;
    22: T504 = 1'h0;
    23: T504 = 1'h0;
    24: T504 = 1'h0;
    25: T504 = 1'h0;
    26: T504 = 1'h0;
    27: T504 = 1'h0;
    28: T504 = 1'h0;
    29: T504 = 1'h0;
    30: T504 = 1'h0;
    31: T504 = 1'h0;
    32: T504 = 1'h0;
    33: T504 = 1'h0;
    34: T504 = 1'h0;
    35: T504 = 1'h0;
    36: T504 = 1'h0;
    37: T504 = 1'h0;
    38: T504 = 1'h0;
    39: T504 = 1'h0;
    40: T504 = 1'h0;
    41: T504 = 1'h0;
    42: T504 = 1'h0;
    43: T504 = 1'h0;
    44: T504 = 1'h0;
    45: T504 = 1'h0;
    46: T504 = 1'h0;
    47: T504 = 1'h0;
    48: T504 = 1'h0;
    49: T504 = 1'h0;
    50: T504 = 1'h0;
    51: T504 = 1'h0;
    52: T504 = 1'h0;
    53: T504 = 1'h0;
    54: T504 = 1'h0;
    55: T504 = 1'h0;
    56: T504 = 1'h0;
    57: T504 = 1'h0;
    58: T504 = 1'h0;
    59: T504 = 1'h0;
    60: T504 = 1'h0;
    61: T504 = 1'h0;
    62: T504 = 1'h0;
    63: T504 = 1'h0;
    64: T504 = 1'h0;
    65: T504 = 1'h0;
    66: T504 = 1'h0;
    67: T504 = 1'h0;
    68: T504 = 1'h0;
    69: T504 = 1'h0;
    70: T504 = 1'h0;
    71: T504 = 1'h0;
    72: T504 = 1'h0;
    73: T504 = 1'h0;
    74: T504 = 1'h0;
    75: T504 = 1'h0;
    76: T504 = 1'h0;
    77: T504 = 1'h0;
    78: T504 = 1'h0;
    79: T504 = 1'h0;
    80: T504 = 1'h0;
    81: T504 = 1'h0;
    82: T504 = 1'h0;
    83: T504 = 1'h0;
    84: T504 = 1'h0;
    85: T504 = 1'h0;
    86: T504 = 1'h0;
    87: T504 = 1'h0;
    88: T504 = 1'h0;
    89: T504 = 1'h0;
    90: T504 = 1'h0;
    91: T504 = 1'h0;
    92: T504 = 1'h0;
    93: T504 = 1'h0;
    94: T504 = 1'h0;
    95: T504 = 1'h0;
    96: T504 = 1'h0;
    97: T504 = 1'h0;
    98: T504 = 1'h0;
    99: T504 = 1'h0;
    100: T504 = 1'h0;
    101: T504 = 1'h0;
    102: T504 = 1'h0;
    103: T504 = 1'h0;
    104: T504 = 1'h0;
    105: T504 = 1'h0;
    106: T504 = 1'h0;
    107: T504 = 1'h0;
    108: T504 = 1'h0;
    109: T504 = 1'h0;
    110: T504 = 1'h0;
    111: T504 = 1'h0;
    112: T504 = 1'h0;
    113: T504 = 1'h0;
    114: T504 = 1'h0;
    115: T504 = 1'h0;
    116: T504 = 1'h0;
    117: T504 = 1'h0;
    118: T504 = 1'h0;
    119: T504 = 1'h0;
    120: T504 = 1'h0;
    121: T504 = 1'h0;
    122: T504 = 1'h0;
    123: T504 = 1'h0;
    124: T504 = 1'h0;
    125: T504 = 1'h0;
    126: T504 = 1'h0;
    127: T504 = 1'h0;
    128: T504 = 1'h0;
    129: T504 = 1'h0;
    130: T504 = 1'h0;
    131: T504 = 1'h0;
    132: T504 = 1'h0;
    133: T504 = 1'h0;
    134: T504 = 1'h0;
    135: T504 = 1'h0;
    136: T504 = 1'h0;
    137: T504 = 1'h0;
    138: T504 = 1'h0;
    139: T504 = 1'h0;
    140: T504 = 1'h0;
    141: T504 = 1'h0;
    142: T504 = 1'h0;
    143: T504 = 1'h0;
    144: T504 = 1'h0;
    145: T504 = 1'h0;
    146: T504 = 1'h0;
    147: T504 = 1'h0;
    148: T504 = 1'h0;
    149: T504 = 1'h0;
    150: T504 = 1'h0;
    151: T504 = 1'h0;
    152: T504 = 1'h0;
    153: T504 = 1'h0;
    154: T504 = 1'h0;
    155: T504 = 1'h0;
    156: T504 = 1'h0;
    157: T504 = 1'h0;
    158: T504 = 1'h0;
    159: T504 = 1'h0;
    160: T504 = 1'h0;
    161: T504 = 1'h0;
    162: T504 = 1'h0;
    163: T504 = 1'h0;
    164: T504 = 1'h0;
    165: T504 = 1'h0;
    166: T504 = 1'h0;
    167: T504 = 1'h0;
    168: T504 = 1'h0;
    169: T504 = 1'h0;
    170: T504 = 1'h0;
    171: T504 = 1'h0;
    172: T504 = 1'h0;
    173: T504 = 1'h0;
    174: T504 = 1'h0;
    175: T504 = 1'h0;
    176: T504 = 1'h0;
    177: T504 = 1'h0;
    178: T504 = 1'h0;
    179: T504 = 1'h0;
    180: T504 = 1'h0;
    181: T504 = 1'h0;
    182: T504 = 1'h0;
    183: T504 = 1'h0;
    184: T504 = 1'h0;
    185: T504 = 1'h0;
    186: T504 = 1'h0;
    187: T504 = 1'h0;
    188: T504 = 1'h0;
    189: T504 = 1'h0;
    190: T504 = 1'h0;
    191: T504 = 1'h0;
    192: T504 = 1'h1;
    193: T504 = 1'h0;
    194: T504 = 1'h0;
    195: T504 = 1'h0;
    196: T504 = 1'h0;
    197: T504 = 1'h0;
    198: T504 = 1'h0;
    199: T504 = 1'h0;
    200: T504 = 1'h0;
    201: T504 = 1'h0;
    202: T504 = 1'h0;
    203: T504 = 1'h0;
    204: T504 = 1'h0;
    205: T504 = 1'h0;
    206: T504 = 1'h0;
    207: T504 = 1'h0;
    208: T504 = 1'h0;
    209: T504 = 1'h0;
    210: T504 = 1'h0;
    211: T504 = 1'h0;
    212: T504 = 1'h0;
    213: T504 = 1'h0;
    214: T504 = 1'h0;
    215: T504 = 1'h0;
    216: T504 = 1'h0;
    217: T504 = 1'h0;
    218: T504 = 1'h0;
    219: T504 = 1'h0;
    220: T504 = 1'h0;
    221: T504 = 1'h0;
    222: T504 = 1'h0;
    223: T504 = 1'h0;
    224: T504 = 1'h0;
    225: T504 = 1'h0;
    226: T504 = 1'h0;
    227: T504 = 1'h0;
    228: T504 = 1'h0;
    229: T504 = 1'h0;
    230: T504 = 1'h0;
    231: T504 = 1'h0;
    232: T504 = 1'h0;
    233: T504 = 1'h0;
    234: T504 = 1'h0;
    235: T504 = 1'h0;
    236: T504 = 1'h0;
    237: T504 = 1'h0;
    238: T504 = 1'h0;
    239: T504 = 1'h0;
    240: T504 = 1'h0;
    241: T504 = 1'h0;
    242: T504 = 1'h0;
    243: T504 = 1'h0;
    244: T504 = 1'h0;
    245: T504 = 1'h0;
    246: T504 = 1'h0;
    247: T504 = 1'h0;
    248: T504 = 1'h0;
    249: T504 = 1'h0;
    250: T504 = 1'h0;
    251: T504 = 1'h0;
    252: T504 = 1'h0;
    253: T504 = 1'h0;
    254: T504 = 1'h0;
    255: T504 = 1'h0;
    256: T504 = 1'h0;
    257: T504 = 1'h0;
    258: T504 = 1'h0;
    259: T504 = 1'h0;
    260: T504 = 1'h0;
    261: T504 = 1'h0;
    262: T504 = 1'h0;
    263: T504 = 1'h0;
    264: T504 = 1'h0;
    265: T504 = 1'h0;
    266: T504 = 1'h0;
    267: T504 = 1'h0;
    268: T504 = 1'h0;
    269: T504 = 1'h0;
    270: T504 = 1'h0;
    271: T504 = 1'h0;
    272: T504 = 1'h0;
    273: T504 = 1'h0;
    274: T504 = 1'h0;
    275: T504 = 1'h0;
    276: T504 = 1'h0;
    277: T504 = 1'h0;
    278: T504 = 1'h0;
    279: T504 = 1'h0;
    280: T504 = 1'h0;
    281: T504 = 1'h0;
    282: T504 = 1'h0;
    283: T504 = 1'h0;
    284: T504 = 1'h0;
    285: T504 = 1'h0;
    286: T504 = 1'h0;
    287: T504 = 1'h0;
    288: T504 = 1'h0;
    289: T504 = 1'h0;
    290: T504 = 1'h0;
    291: T504 = 1'h0;
    292: T504 = 1'h0;
    293: T504 = 1'h0;
    294: T504 = 1'h0;
    295: T504 = 1'h0;
    296: T504 = 1'h0;
    297: T504 = 1'h0;
    298: T504 = 1'h0;
    299: T504 = 1'h0;
    300: T504 = 1'h0;
    301: T504 = 1'h0;
    302: T504 = 1'h0;
    303: T504 = 1'h0;
    304: T504 = 1'h0;
    305: T504 = 1'h0;
    306: T504 = 1'h0;
    307: T504 = 1'h0;
    308: T504 = 1'h0;
    309: T504 = 1'h0;
    310: T504 = 1'h0;
    311: T504 = 1'h0;
    312: T504 = 1'h0;
    313: T504 = 1'h0;
    314: T504 = 1'h0;
    315: T504 = 1'h0;
    316: T504 = 1'h0;
    317: T504 = 1'h0;
    318: T504 = 1'h0;
    319: T504 = 1'h0;
    320: T504 = 1'h0;
    321: T504 = 1'h0;
    322: T504 = 1'h0;
    323: T504 = 1'h0;
    324: T504 = 1'h0;
    325: T504 = 1'h0;
    326: T504 = 1'h0;
    327: T504 = 1'h0;
    328: T504 = 1'h0;
    329: T504 = 1'h0;
    330: T504 = 1'h0;
    331: T504 = 1'h0;
    332: T504 = 1'h0;
    333: T504 = 1'h0;
    334: T504 = 1'h0;
    335: T504 = 1'h0;
    336: T504 = 1'h0;
    337: T504 = 1'h0;
    338: T504 = 1'h0;
    339: T504 = 1'h0;
    340: T504 = 1'h0;
    341: T504 = 1'h0;
    342: T504 = 1'h0;
    343: T504 = 1'h0;
    344: T504 = 1'h0;
    345: T504 = 1'h0;
    346: T504 = 1'h0;
    347: T504 = 1'h0;
    348: T504 = 1'h0;
    349: T504 = 1'h0;
    350: T504 = 1'h0;
    351: T504 = 1'h0;
    352: T504 = 1'h0;
    353: T504 = 1'h0;
    354: T504 = 1'h0;
    355: T504 = 1'h0;
    356: T504 = 1'h0;
    357: T504 = 1'h0;
    358: T504 = 1'h0;
    359: T504 = 1'h0;
    360: T504 = 1'h0;
    361: T504 = 1'h0;
    362: T504 = 1'h0;
    363: T504 = 1'h0;
    364: T504 = 1'h0;
    365: T504 = 1'h0;
    366: T504 = 1'h0;
    367: T504 = 1'h0;
    368: T504 = 1'h0;
    369: T504 = 1'h0;
    370: T504 = 1'h0;
    371: T504 = 1'h0;
    372: T504 = 1'h0;
    373: T504 = 1'h0;
    374: T504 = 1'h0;
    375: T504 = 1'h0;
    376: T504 = 1'h0;
    377: T504 = 1'h0;
    378: T504 = 1'h0;
    379: T504 = 1'h0;
    380: T504 = 1'h0;
    381: T504 = 1'h0;
    382: T504 = 1'h0;
    383: T504 = 1'h0;
    384: T504 = 1'h0;
    385: T504 = 1'h0;
    386: T504 = 1'h0;
    387: T504 = 1'h0;
    388: T504 = 1'h0;
    389: T504 = 1'h0;
    390: T504 = 1'h0;
    391: T504 = 1'h0;
    392: T504 = 1'h0;
    393: T504 = 1'h0;
    394: T504 = 1'h0;
    395: T504 = 1'h0;
    396: T504 = 1'h0;
    397: T504 = 1'h0;
    398: T504 = 1'h0;
    399: T504 = 1'h0;
    400: T504 = 1'h0;
    401: T504 = 1'h0;
    402: T504 = 1'h0;
    403: T504 = 1'h0;
    404: T504 = 1'h0;
    405: T504 = 1'h0;
    406: T504 = 1'h0;
    407: T504 = 1'h0;
    408: T504 = 1'h0;
    409: T504 = 1'h0;
    410: T504 = 1'h0;
    411: T504 = 1'h0;
    412: T504 = 1'h0;
    413: T504 = 1'h0;
    414: T504 = 1'h0;
    415: T504 = 1'h0;
    416: T504 = 1'h0;
    417: T504 = 1'h0;
    418: T504 = 1'h0;
    419: T504 = 1'h0;
    420: T504 = 1'h0;
    421: T504 = 1'h0;
    422: T504 = 1'h0;
    423: T504 = 1'h0;
    424: T504 = 1'h0;
    425: T504 = 1'h0;
    426: T504 = 1'h0;
    427: T504 = 1'h0;
    428: T504 = 1'h0;
    429: T504 = 1'h0;
    430: T504 = 1'h0;
    431: T504 = 1'h0;
    432: T504 = 1'h0;
    433: T504 = 1'h0;
    434: T504 = 1'h0;
    435: T504 = 1'h0;
    436: T504 = 1'h0;
    437: T504 = 1'h0;
    438: T504 = 1'h0;
    439: T504 = 1'h0;
    440: T504 = 1'h0;
    441: T504 = 1'h0;
    442: T504 = 1'h0;
    443: T504 = 1'h0;
    444: T504 = 1'h0;
    445: T504 = 1'h0;
    446: T504 = 1'h0;
    447: T504 = 1'h0;
    448: T504 = 1'h0;
    449: T504 = 1'h0;
    450: T504 = 1'h0;
    451: T504 = 1'h0;
    452: T504 = 1'h0;
    453: T504 = 1'h0;
    454: T504 = 1'h0;
    455: T504 = 1'h0;
    456: T504 = 1'h0;
    457: T504 = 1'h0;
    458: T504 = 1'h0;
    459: T504 = 1'h0;
    460: T504 = 1'h0;
    461: T504 = 1'h0;
    462: T504 = 1'h0;
    463: T504 = 1'h0;
    464: T504 = 1'h0;
    465: T504 = 1'h0;
    466: T504 = 1'h0;
    467: T504 = 1'h0;
    468: T504 = 1'h0;
    469: T504 = 1'h0;
    470: T504 = 1'h0;
    471: T504 = 1'h0;
    472: T504 = 1'h0;
    473: T504 = 1'h0;
    474: T504 = 1'h0;
    475: T504 = 1'h0;
    476: T504 = 1'h0;
    477: T504 = 1'h0;
    478: T504 = 1'h0;
    479: T504 = 1'h0;
    480: T504 = 1'h0;
    481: T504 = 1'h0;
    482: T504 = 1'h0;
    483: T504 = 1'h0;
    484: T504 = 1'h0;
    485: T504 = 1'h0;
    486: T504 = 1'h0;
    487: T504 = 1'h0;
    488: T504 = 1'h0;
    489: T504 = 1'h0;
    490: T504 = 1'h0;
    491: T504 = 1'h0;
    492: T504 = 1'h0;
    493: T504 = 1'h0;
    494: T504 = 1'h0;
    495: T504 = 1'h0;
    496: T504 = 1'h0;
    497: T504 = 1'h0;
    498: T504 = 1'h0;
    499: T504 = 1'h0;
    500: T504 = 1'h0;
    501: T504 = 1'h0;
    502: T504 = 1'h0;
    503: T504 = 1'h0;
    504: T504 = 1'h0;
    505: T504 = 1'h0;
    506: T504 = 1'h0;
    507: T504 = 1'h0;
    508: T504 = 1'h0;
    509: T504 = 1'h0;
    510: T504 = 1'h0;
    511: T504 = 1'h0;
    512: T504 = 1'h0;
    513: T504 = 1'h0;
    514: T504 = 1'h0;
    515: T504 = 1'h0;
    516: T504 = 1'h0;
    517: T504 = 1'h0;
    518: T504 = 1'h0;
    519: T504 = 1'h0;
    520: T504 = 1'h0;
    521: T504 = 1'h0;
    522: T504 = 1'h0;
    523: T504 = 1'h0;
    524: T504 = 1'h0;
    525: T504 = 1'h0;
    526: T504 = 1'h0;
    527: T504 = 1'h0;
    528: T504 = 1'h0;
    529: T504 = 1'h0;
    530: T504 = 1'h0;
    531: T504 = 1'h0;
    532: T504 = 1'h0;
    533: T504 = 1'h0;
    534: T504 = 1'h0;
    535: T504 = 1'h0;
    536: T504 = 1'h0;
    537: T504 = 1'h0;
    538: T504 = 1'h0;
    539: T504 = 1'h0;
    540: T504 = 1'h0;
    541: T504 = 1'h0;
    542: T504 = 1'h0;
    543: T504 = 1'h0;
    544: T504 = 1'h0;
    545: T504 = 1'h0;
    546: T504 = 1'h0;
    547: T504 = 1'h0;
    548: T504 = 1'h0;
    549: T504 = 1'h0;
    550: T504 = 1'h0;
    551: T504 = 1'h0;
    552: T504 = 1'h0;
    553: T504 = 1'h0;
    554: T504 = 1'h0;
    555: T504 = 1'h0;
    556: T504 = 1'h0;
    557: T504 = 1'h0;
    558: T504 = 1'h0;
    559: T504 = 1'h0;
    560: T504 = 1'h0;
    561: T504 = 1'h0;
    562: T504 = 1'h0;
    563: T504 = 1'h0;
    564: T504 = 1'h0;
    565: T504 = 1'h0;
    566: T504 = 1'h0;
    567: T504 = 1'h0;
    568: T504 = 1'h0;
    569: T504 = 1'h0;
    570: T504 = 1'h0;
    571: T504 = 1'h0;
    572: T504 = 1'h0;
    573: T504 = 1'h0;
    574: T504 = 1'h0;
    575: T504 = 1'h0;
    576: T504 = 1'h0;
    577: T504 = 1'h0;
    578: T504 = 1'h0;
    579: T504 = 1'h0;
    580: T504 = 1'h0;
    581: T504 = 1'h0;
    582: T504 = 1'h0;
    583: T504 = 1'h0;
    584: T504 = 1'h0;
    585: T504 = 1'h0;
    586: T504 = 1'h0;
    587: T504 = 1'h0;
    588: T504 = 1'h0;
    589: T504 = 1'h0;
    590: T504 = 1'h0;
    591: T504 = 1'h0;
    592: T504 = 1'h0;
    593: T504 = 1'h0;
    594: T504 = 1'h0;
    595: T504 = 1'h0;
    596: T504 = 1'h0;
    597: T504 = 1'h0;
    598: T504 = 1'h0;
    599: T504 = 1'h0;
    600: T504 = 1'h0;
    601: T504 = 1'h0;
    602: T504 = 1'h0;
    603: T504 = 1'h0;
    604: T504 = 1'h0;
    605: T504 = 1'h0;
    606: T504 = 1'h0;
    607: T504 = 1'h0;
    608: T504 = 1'h0;
    609: T504 = 1'h0;
    610: T504 = 1'h0;
    611: T504 = 1'h0;
    612: T504 = 1'h0;
    613: T504 = 1'h0;
    614: T504 = 1'h0;
    615: T504 = 1'h0;
    616: T504 = 1'h0;
    617: T504 = 1'h0;
    618: T504 = 1'h0;
    619: T504 = 1'h0;
    620: T504 = 1'h0;
    621: T504 = 1'h0;
    622: T504 = 1'h0;
    623: T504 = 1'h0;
    624: T504 = 1'h0;
    625: T504 = 1'h0;
    626: T504 = 1'h0;
    627: T504 = 1'h0;
    628: T504 = 1'h0;
    629: T504 = 1'h0;
    630: T504 = 1'h0;
    631: T504 = 1'h0;
    632: T504 = 1'h0;
    633: T504 = 1'h0;
    634: T504 = 1'h0;
    635: T504 = 1'h0;
    636: T504 = 1'h0;
    637: T504 = 1'h0;
    638: T504 = 1'h0;
    639: T504 = 1'h0;
    640: T504 = 1'h0;
    641: T504 = 1'h0;
    642: T504 = 1'h0;
    643: T504 = 1'h0;
    644: T504 = 1'h0;
    645: T504 = 1'h0;
    646: T504 = 1'h0;
    647: T504 = 1'h0;
    648: T504 = 1'h0;
    649: T504 = 1'h0;
    650: T504 = 1'h0;
    651: T504 = 1'h0;
    652: T504 = 1'h0;
    653: T504 = 1'h0;
    654: T504 = 1'h0;
    655: T504 = 1'h0;
    656: T504 = 1'h0;
    657: T504 = 1'h0;
    658: T504 = 1'h0;
    659: T504 = 1'h0;
    660: T504 = 1'h0;
    661: T504 = 1'h0;
    662: T504 = 1'h0;
    663: T504 = 1'h0;
    664: T504 = 1'h0;
    665: T504 = 1'h0;
    666: T504 = 1'h0;
    667: T504 = 1'h0;
    668: T504 = 1'h0;
    669: T504 = 1'h0;
    670: T504 = 1'h0;
    671: T504 = 1'h0;
    672: T504 = 1'h0;
    673: T504 = 1'h0;
    674: T504 = 1'h0;
    675: T504 = 1'h0;
    676: T504 = 1'h0;
    677: T504 = 1'h0;
    678: T504 = 1'h0;
    679: T504 = 1'h0;
    680: T504 = 1'h0;
    681: T504 = 1'h0;
    682: T504 = 1'h0;
    683: T504 = 1'h0;
    684: T504 = 1'h0;
    685: T504 = 1'h0;
    686: T504 = 1'h0;
    687: T504 = 1'h0;
    688: T504 = 1'h0;
    689: T504 = 1'h0;
    690: T504 = 1'h0;
    691: T504 = 1'h0;
    692: T504 = 1'h0;
    693: T504 = 1'h0;
    694: T504 = 1'h0;
    695: T504 = 1'h0;
    696: T504 = 1'h0;
    697: T504 = 1'h0;
    698: T504 = 1'h0;
    699: T504 = 1'h0;
    700: T504 = 1'h0;
    701: T504 = 1'h0;
    702: T504 = 1'h0;
    703: T504 = 1'h0;
    704: T504 = 1'h0;
    705: T504 = 1'h0;
    706: T504 = 1'h0;
    707: T504 = 1'h0;
    708: T504 = 1'h0;
    709: T504 = 1'h0;
    710: T504 = 1'h0;
    711: T504 = 1'h0;
    712: T504 = 1'h0;
    713: T504 = 1'h0;
    714: T504 = 1'h0;
    715: T504 = 1'h0;
    716: T504 = 1'h0;
    717: T504 = 1'h0;
    718: T504 = 1'h0;
    719: T504 = 1'h0;
    720: T504 = 1'h0;
    721: T504 = 1'h0;
    722: T504 = 1'h0;
    723: T504 = 1'h0;
    724: T504 = 1'h0;
    725: T504 = 1'h0;
    726: T504 = 1'h0;
    727: T504 = 1'h0;
    728: T504 = 1'h0;
    729: T504 = 1'h0;
    730: T504 = 1'h0;
    731: T504 = 1'h0;
    732: T504 = 1'h0;
    733: T504 = 1'h0;
    734: T504 = 1'h0;
    735: T504 = 1'h0;
    736: T504 = 1'h0;
    737: T504 = 1'h0;
    738: T504 = 1'h0;
    739: T504 = 1'h0;
    740: T504 = 1'h0;
    741: T504 = 1'h0;
    742: T504 = 1'h0;
    743: T504 = 1'h0;
    744: T504 = 1'h0;
    745: T504 = 1'h0;
    746: T504 = 1'h0;
    747: T504 = 1'h0;
    748: T504 = 1'h0;
    749: T504 = 1'h0;
    750: T504 = 1'h0;
    751: T504 = 1'h0;
    752: T504 = 1'h0;
    753: T504 = 1'h0;
    754: T504 = 1'h0;
    755: T504 = 1'h0;
    756: T504 = 1'h0;
    757: T504 = 1'h0;
    758: T504 = 1'h0;
    759: T504 = 1'h0;
    760: T504 = 1'h0;
    761: T504 = 1'h0;
    762: T504 = 1'h0;
    763: T504 = 1'h0;
    764: T504 = 1'h0;
    765: T504 = 1'h0;
    766: T504 = 1'h0;
    767: T504 = 1'h0;
    768: T504 = 1'h0;
    769: T504 = 1'h0;
    770: T504 = 1'h0;
    771: T504 = 1'h0;
    772: T504 = 1'h0;
    773: T504 = 1'h0;
    774: T504 = 1'h0;
    775: T504 = 1'h0;
    776: T504 = 1'h0;
    777: T504 = 1'h0;
    778: T504 = 1'h0;
    779: T504 = 1'h0;
    780: T504 = 1'h0;
    781: T504 = 1'h0;
    782: T504 = 1'h0;
    783: T504 = 1'h0;
    784: T504 = 1'h0;
    785: T504 = 1'h0;
    786: T504 = 1'h0;
    787: T504 = 1'h0;
    788: T504 = 1'h0;
    789: T504 = 1'h0;
    790: T504 = 1'h0;
    791: T504 = 1'h0;
    792: T504 = 1'h0;
    793: T504 = 1'h0;
    794: T504 = 1'h0;
    795: T504 = 1'h0;
    796: T504 = 1'h0;
    797: T504 = 1'h0;
    798: T504 = 1'h0;
    799: T504 = 1'h0;
    800: T504 = 1'h0;
    801: T504 = 1'h0;
    802: T504 = 1'h0;
    803: T504 = 1'h0;
    804: T504 = 1'h0;
    805: T504 = 1'h0;
    806: T504 = 1'h0;
    807: T504 = 1'h0;
    808: T504 = 1'h0;
    809: T504 = 1'h0;
    810: T504 = 1'h0;
    811: T504 = 1'h0;
    812: T504 = 1'h0;
    813: T504 = 1'h0;
    814: T504 = 1'h0;
    815: T504 = 1'h0;
    816: T504 = 1'h0;
    817: T504 = 1'h0;
    818: T504 = 1'h0;
    819: T504 = 1'h0;
    820: T504 = 1'h0;
    821: T504 = 1'h0;
    822: T504 = 1'h0;
    823: T504 = 1'h0;
    824: T504 = 1'h0;
    825: T504 = 1'h0;
    826: T504 = 1'h0;
    827: T504 = 1'h0;
    828: T504 = 1'h0;
    829: T504 = 1'h0;
    830: T504 = 1'h0;
    831: T504 = 1'h0;
    832: T504 = 1'h0;
    833: T504 = 1'h0;
    834: T504 = 1'h0;
    835: T504 = 1'h0;
    836: T504 = 1'h0;
    837: T504 = 1'h0;
    838: T504 = 1'h0;
    839: T504 = 1'h0;
    840: T504 = 1'h0;
    841: T504 = 1'h0;
    842: T504 = 1'h0;
    843: T504 = 1'h0;
    844: T504 = 1'h0;
    845: T504 = 1'h0;
    846: T504 = 1'h0;
    847: T504 = 1'h0;
    848: T504 = 1'h0;
    849: T504 = 1'h0;
    850: T504 = 1'h0;
    851: T504 = 1'h0;
    852: T504 = 1'h0;
    853: T504 = 1'h0;
    854: T504 = 1'h0;
    855: T504 = 1'h0;
    856: T504 = 1'h0;
    857: T504 = 1'h0;
    858: T504 = 1'h0;
    859: T504 = 1'h0;
    860: T504 = 1'h0;
    861: T504 = 1'h0;
    862: T504 = 1'h0;
    863: T504 = 1'h0;
    864: T504 = 1'h0;
    865: T504 = 1'h0;
    866: T504 = 1'h0;
    867: T504 = 1'h0;
    868: T504 = 1'h0;
    869: T504 = 1'h0;
    870: T504 = 1'h0;
    871: T504 = 1'h0;
    872: T504 = 1'h0;
    873: T504 = 1'h0;
    874: T504 = 1'h0;
    875: T504 = 1'h0;
    876: T504 = 1'h0;
    877: T504 = 1'h0;
    878: T504 = 1'h0;
    879: T504 = 1'h0;
    880: T504 = 1'h0;
    881: T504 = 1'h0;
    882: T504 = 1'h0;
    883: T504 = 1'h0;
    884: T504 = 1'h0;
    885: T504 = 1'h0;
    886: T504 = 1'h0;
    887: T504 = 1'h0;
    888: T504 = 1'h0;
    889: T504 = 1'h0;
    890: T504 = 1'h0;
    891: T504 = 1'h0;
    892: T504 = 1'h0;
    893: T504 = 1'h0;
    894: T504 = 1'h0;
    895: T504 = 1'h0;
    896: T504 = 1'h0;
    897: T504 = 1'h0;
    898: T504 = 1'h0;
    899: T504 = 1'h0;
    900: T504 = 1'h0;
    901: T504 = 1'h0;
    902: T504 = 1'h0;
    903: T504 = 1'h0;
    904: T504 = 1'h0;
    905: T504 = 1'h0;
    906: T504 = 1'h0;
    907: T504 = 1'h0;
    908: T504 = 1'h0;
    909: T504 = 1'h0;
    910: T504 = 1'h0;
    911: T504 = 1'h0;
    912: T504 = 1'h0;
    913: T504 = 1'h0;
    914: T504 = 1'h0;
    915: T504 = 1'h0;
    916: T504 = 1'h0;
    917: T504 = 1'h0;
    918: T504 = 1'h0;
    919: T504 = 1'h0;
    920: T504 = 1'h0;
    921: T504 = 1'h0;
    922: T504 = 1'h0;
    923: T504 = 1'h0;
    924: T504 = 1'h0;
    925: T504 = 1'h0;
    926: T504 = 1'h0;
    927: T504 = 1'h0;
    928: T504 = 1'h0;
    929: T504 = 1'h0;
    930: T504 = 1'h0;
    931: T504 = 1'h0;
    932: T504 = 1'h0;
    933: T504 = 1'h0;
    934: T504 = 1'h0;
    935: T504 = 1'h0;
    936: T504 = 1'h0;
    937: T504 = 1'h0;
    938: T504 = 1'h0;
    939: T504 = 1'h0;
    940: T504 = 1'h0;
    941: T504 = 1'h0;
    942: T504 = 1'h0;
    943: T504 = 1'h0;
    944: T504 = 1'h0;
    945: T504 = 1'h0;
    946: T504 = 1'h0;
    947: T504 = 1'h0;
    948: T504 = 1'h0;
    949: T504 = 1'h0;
    950: T504 = 1'h0;
    951: T504 = 1'h0;
    952: T504 = 1'h0;
    953: T504 = 1'h0;
    954: T504 = 1'h0;
    955: T504 = 1'h0;
    956: T504 = 1'h0;
    957: T504 = 1'h0;
    958: T504 = 1'h0;
    959: T504 = 1'h0;
    960: T504 = 1'h0;
    961: T504 = 1'h0;
    962: T504 = 1'h0;
    963: T504 = 1'h0;
    964: T504 = 1'h0;
    965: T504 = 1'h0;
    966: T504 = 1'h0;
    967: T504 = 1'h0;
    968: T504 = 1'h0;
    969: T504 = 1'h0;
    970: T504 = 1'h0;
    971: T504 = 1'h0;
    972: T504 = 1'h0;
    973: T504 = 1'h0;
    974: T504 = 1'h0;
    975: T504 = 1'h0;
    976: T504 = 1'h0;
    977: T504 = 1'h0;
    978: T504 = 1'h0;
    979: T504 = 1'h0;
    980: T504 = 1'h0;
    981: T504 = 1'h0;
    982: T504 = 1'h0;
    983: T504 = 1'h0;
    984: T504 = 1'h0;
    985: T504 = 1'h0;
    986: T504 = 1'h0;
    987: T504 = 1'h0;
    988: T504 = 1'h0;
    989: T504 = 1'h0;
    990: T504 = 1'h0;
    991: T504 = 1'h0;
    992: T504 = 1'h0;
    993: T504 = 1'h0;
    994: T504 = 1'h0;
    995: T504 = 1'h0;
    996: T504 = 1'h0;
    997: T504 = 1'h0;
    998: T504 = 1'h0;
    999: T504 = 1'h0;
    1000: T504 = 1'h0;
    1001: T504 = 1'h0;
    1002: T504 = 1'h0;
    1003: T504 = 1'h0;
    1004: T504 = 1'h0;
    1005: T504 = 1'h0;
    1006: T504 = 1'h0;
    1007: T504 = 1'h0;
    1008: T504 = 1'h0;
    1009: T504 = 1'h0;
    1010: T504 = 1'h0;
    1011: T504 = 1'h0;
    1012: T504 = 1'h0;
    1013: T504 = 1'h0;
    1014: T504 = 1'h0;
    1015: T504 = 1'h0;
    1016: T504 = 1'h0;
    1017: T504 = 1'h0;
    1018: T504 = 1'h0;
    1019: T504 = 1'h0;
    1020: T504 = 1'h0;
    1021: T504 = 1'h0;
    1022: T504 = 1'h0;
    1023: T504 = 1'h0;
    1024: T504 = 1'h0;
    1025: T504 = 1'h0;
    1026: T504 = 1'h0;
    1027: T504 = 1'h0;
    1028: T504 = 1'h0;
    1029: T504 = 1'h0;
    1030: T504 = 1'h0;
    1031: T504 = 1'h0;
    1032: T504 = 1'h0;
    1033: T504 = 1'h0;
    1034: T504 = 1'h0;
    1035: T504 = 1'h0;
    1036: T504 = 1'h0;
    1037: T504 = 1'h0;
    1038: T504 = 1'h0;
    1039: T504 = 1'h0;
    1040: T504 = 1'h0;
    1041: T504 = 1'h0;
    1042: T504 = 1'h0;
    1043: T504 = 1'h0;
    1044: T504 = 1'h0;
    1045: T504 = 1'h0;
    1046: T504 = 1'h0;
    1047: T504 = 1'h0;
    1048: T504 = 1'h0;
    1049: T504 = 1'h0;
    1050: T504 = 1'h0;
    1051: T504 = 1'h0;
    1052: T504 = 1'h0;
    1053: T504 = 1'h0;
    1054: T504 = 1'h0;
    1055: T504 = 1'h0;
    1056: T504 = 1'h0;
    1057: T504 = 1'h0;
    1058: T504 = 1'h0;
    1059: T504 = 1'h0;
    1060: T504 = 1'h0;
    1061: T504 = 1'h0;
    1062: T504 = 1'h0;
    1063: T504 = 1'h0;
    1064: T504 = 1'h0;
    1065: T504 = 1'h0;
    1066: T504 = 1'h0;
    1067: T504 = 1'h0;
    1068: T504 = 1'h0;
    1069: T504 = 1'h0;
    1070: T504 = 1'h0;
    1071: T504 = 1'h0;
    1072: T504 = 1'h0;
    1073: T504 = 1'h0;
    1074: T504 = 1'h0;
    1075: T504 = 1'h0;
    1076: T504 = 1'h0;
    1077: T504 = 1'h0;
    1078: T504 = 1'h0;
    1079: T504 = 1'h0;
    1080: T504 = 1'h0;
    1081: T504 = 1'h0;
    1082: T504 = 1'h0;
    1083: T504 = 1'h0;
    1084: T504 = 1'h0;
    1085: T504 = 1'h0;
    1086: T504 = 1'h0;
    1087: T504 = 1'h0;
    1088: T504 = 1'h0;
    1089: T504 = 1'h0;
    1090: T504 = 1'h0;
    1091: T504 = 1'h0;
    1092: T504 = 1'h0;
    1093: T504 = 1'h0;
    1094: T504 = 1'h0;
    1095: T504 = 1'h0;
    1096: T504 = 1'h0;
    1097: T504 = 1'h0;
    1098: T504 = 1'h0;
    1099: T504 = 1'h0;
    1100: T504 = 1'h0;
    1101: T504 = 1'h0;
    1102: T504 = 1'h0;
    1103: T504 = 1'h0;
    1104: T504 = 1'h0;
    1105: T504 = 1'h0;
    1106: T504 = 1'h0;
    1107: T504 = 1'h0;
    1108: T504 = 1'h0;
    1109: T504 = 1'h0;
    1110: T504 = 1'h0;
    1111: T504 = 1'h0;
    1112: T504 = 1'h0;
    1113: T504 = 1'h0;
    1114: T504 = 1'h0;
    1115: T504 = 1'h0;
    1116: T504 = 1'h0;
    1117: T504 = 1'h0;
    1118: T504 = 1'h0;
    1119: T504 = 1'h0;
    1120: T504 = 1'h0;
    1121: T504 = 1'h0;
    1122: T504 = 1'h0;
    1123: T504 = 1'h0;
    1124: T504 = 1'h0;
    1125: T504 = 1'h0;
    1126: T504 = 1'h0;
    1127: T504 = 1'h0;
    1128: T504 = 1'h0;
    1129: T504 = 1'h0;
    1130: T504 = 1'h0;
    1131: T504 = 1'h0;
    1132: T504 = 1'h0;
    1133: T504 = 1'h0;
    1134: T504 = 1'h0;
    1135: T504 = 1'h0;
    1136: T504 = 1'h0;
    1137: T504 = 1'h0;
    1138: T504 = 1'h0;
    1139: T504 = 1'h0;
    1140: T504 = 1'h0;
    1141: T504 = 1'h0;
    1142: T504 = 1'h0;
    1143: T504 = 1'h0;
    1144: T504 = 1'h0;
    1145: T504 = 1'h0;
    1146: T504 = 1'h0;
    1147: T504 = 1'h0;
    1148: T504 = 1'h0;
    1149: T504 = 1'h0;
    1150: T504 = 1'h0;
    1151: T504 = 1'h0;
    1152: T504 = 1'h0;
    1153: T504 = 1'h0;
    1154: T504 = 1'h0;
    1155: T504 = 1'h0;
    1156: T504 = 1'h0;
    1157: T504 = 1'h0;
    1158: T504 = 1'h0;
    1159: T504 = 1'h0;
    1160: T504 = 1'h0;
    1161: T504 = 1'h0;
    1162: T504 = 1'h0;
    1163: T504 = 1'h0;
    1164: T504 = 1'h0;
    1165: T504 = 1'h0;
    1166: T504 = 1'h0;
    1167: T504 = 1'h0;
    1168: T504 = 1'h0;
    1169: T504 = 1'h0;
    1170: T504 = 1'h0;
    1171: T504 = 1'h0;
    1172: T504 = 1'h0;
    1173: T504 = 1'h0;
    1174: T504 = 1'h0;
    1175: T504 = 1'h0;
    1176: T504 = 1'h0;
    1177: T504 = 1'h0;
    1178: T504 = 1'h0;
    1179: T504 = 1'h0;
    1180: T504 = 1'h0;
    1181: T504 = 1'h0;
    1182: T504 = 1'h0;
    1183: T504 = 1'h0;
    1184: T504 = 1'h0;
    1185: T504 = 1'h0;
    1186: T504 = 1'h0;
    1187: T504 = 1'h0;
    1188: T504 = 1'h0;
    1189: T504 = 1'h0;
    1190: T504 = 1'h0;
    1191: T504 = 1'h0;
    1192: T504 = 1'h0;
    1193: T504 = 1'h0;
    1194: T504 = 1'h0;
    1195: T504 = 1'h0;
    1196: T504 = 1'h0;
    1197: T504 = 1'h0;
    1198: T504 = 1'h0;
    1199: T504 = 1'h0;
    1200: T504 = 1'h0;
    1201: T504 = 1'h0;
    1202: T504 = 1'h0;
    1203: T504 = 1'h0;
    1204: T504 = 1'h0;
    1205: T504 = 1'h0;
    1206: T504 = 1'h0;
    1207: T504 = 1'h0;
    1208: T504 = 1'h0;
    1209: T504 = 1'h0;
    1210: T504 = 1'h0;
    1211: T504 = 1'h0;
    1212: T504 = 1'h0;
    1213: T504 = 1'h0;
    1214: T504 = 1'h0;
    1215: T504 = 1'h0;
    1216: T504 = 1'h0;
    1217: T504 = 1'h0;
    1218: T504 = 1'h0;
    1219: T504 = 1'h0;
    1220: T504 = 1'h0;
    1221: T504 = 1'h0;
    1222: T504 = 1'h0;
    1223: T504 = 1'h0;
    1224: T504 = 1'h0;
    1225: T504 = 1'h0;
    1226: T504 = 1'h0;
    1227: T504 = 1'h0;
    1228: T504 = 1'h0;
    1229: T504 = 1'h0;
    1230: T504 = 1'h0;
    1231: T504 = 1'h0;
    1232: T504 = 1'h0;
    1233: T504 = 1'h0;
    1234: T504 = 1'h0;
    1235: T504 = 1'h0;
    1236: T504 = 1'h0;
    1237: T504 = 1'h0;
    1238: T504 = 1'h0;
    1239: T504 = 1'h0;
    1240: T504 = 1'h0;
    1241: T504 = 1'h0;
    1242: T504 = 1'h0;
    1243: T504 = 1'h0;
    1244: T504 = 1'h0;
    1245: T504 = 1'h0;
    1246: T504 = 1'h0;
    1247: T504 = 1'h0;
    1248: T504 = 1'h0;
    1249: T504 = 1'h0;
    1250: T504 = 1'h0;
    1251: T504 = 1'h0;
    1252: T504 = 1'h0;
    1253: T504 = 1'h0;
    1254: T504 = 1'h0;
    1255: T504 = 1'h0;
    1256: T504 = 1'h0;
    1257: T504 = 1'h0;
    1258: T504 = 1'h0;
    1259: T504 = 1'h0;
    1260: T504 = 1'h0;
    1261: T504 = 1'h0;
    1262: T504 = 1'h0;
    1263: T504 = 1'h0;
    1264: T504 = 1'h0;
    1265: T504 = 1'h0;
    1266: T504 = 1'h0;
    1267: T504 = 1'h0;
    1268: T504 = 1'h0;
    1269: T504 = 1'h0;
    1270: T504 = 1'h0;
    1271: T504 = 1'h0;
    1272: T504 = 1'h0;
    1273: T504 = 1'h0;
    1274: T504 = 1'h0;
    1275: T504 = 1'h0;
    1276: T504 = 1'h0;
    1277: T504 = 1'h0;
    1278: T504 = 1'h0;
    1279: T504 = 1'h0;
    1280: T504 = 1'h1;
    1281: T504 = 1'h1;
    1282: T504 = 1'h1;
    1283: T504 = 1'h1;
    1284: T504 = 1'h1;
    1285: T504 = 1'h1;
    1286: T504 = 1'h1;
    1287: T504 = 1'h1;
    1288: T504 = 1'h1;
    1289: T504 = 1'h1;
    1290: T504 = 1'h1;
    1291: T504 = 1'h1;
    1292: T504 = 1'h1;
    1293: T504 = 1'h1;
    1294: T504 = 1'h1;
    1295: T504 = 1'h1;
    1296: T504 = 1'h0;
    1297: T504 = 1'h0;
    1298: T504 = 1'h0;
    1299: T504 = 1'h0;
    1300: T504 = 1'h0;
    1301: T504 = 1'h0;
    1302: T504 = 1'h0;
    1303: T504 = 1'h0;
    1304: T504 = 1'h0;
    1305: T504 = 1'h0;
    1306: T504 = 1'h0;
    1307: T504 = 1'h0;
    1308: T504 = 1'h0;
    1309: T504 = 1'h1;
    1310: T504 = 1'h1;
    1311: T504 = 1'h1;
    1312: T504 = 1'h1;
    1313: T504 = 1'h0;
    1314: T504 = 1'h0;
    1315: T504 = 1'h0;
    1316: T504 = 1'h0;
    1317: T504 = 1'h0;
    1318: T504 = 1'h0;
    1319: T504 = 1'h0;
    1320: T504 = 1'h0;
    1321: T504 = 1'h0;
    1322: T504 = 1'h0;
    1323: T504 = 1'h0;
    1324: T504 = 1'h0;
    1325: T504 = 1'h0;
    1326: T504 = 1'h0;
    1327: T504 = 1'h0;
    1328: T504 = 1'h0;
    1329: T504 = 1'h0;
    1330: T504 = 1'h0;
    1331: T504 = 1'h0;
    1332: T504 = 1'h0;
    1333: T504 = 1'h0;
    1334: T504 = 1'h0;
    1335: T504 = 1'h0;
    1336: T504 = 1'h0;
    1337: T504 = 1'h0;
    1338: T504 = 1'h0;
    1339: T504 = 1'h0;
    1340: T504 = 1'h0;
    1341: T504 = 1'h0;
    1342: T504 = 1'h0;
    1343: T504 = 1'h0;
    1344: T504 = 1'h0;
    1345: T504 = 1'h0;
    1346: T504 = 1'h0;
    1347: T504 = 1'h0;
    1348: T504 = 1'h0;
    1349: T504 = 1'h0;
    1350: T504 = 1'h0;
    1351: T504 = 1'h0;
    1352: T504 = 1'h0;
    1353: T504 = 1'h0;
    1354: T504 = 1'h0;
    1355: T504 = 1'h0;
    1356: T504 = 1'h0;
    1357: T504 = 1'h0;
    1358: T504 = 1'h0;
    1359: T504 = 1'h0;
    1360: T504 = 1'h0;
    1361: T504 = 1'h0;
    1362: T504 = 1'h0;
    1363: T504 = 1'h0;
    1364: T504 = 1'h0;
    1365: T504 = 1'h0;
    1366: T504 = 1'h0;
    1367: T504 = 1'h0;
    1368: T504 = 1'h0;
    1369: T504 = 1'h0;
    1370: T504 = 1'h0;
    1371: T504 = 1'h0;
    1372: T504 = 1'h0;
    1373: T504 = 1'h0;
    1374: T504 = 1'h0;
    1375: T504 = 1'h0;
    1376: T504 = 1'h0;
    1377: T504 = 1'h0;
    1378: T504 = 1'h0;
    1379: T504 = 1'h0;
    1380: T504 = 1'h0;
    1381: T504 = 1'h0;
    1382: T504 = 1'h0;
    1383: T504 = 1'h0;
    1384: T504 = 1'h0;
    1385: T504 = 1'h0;
    1386: T504 = 1'h0;
    1387: T504 = 1'h0;
    1388: T504 = 1'h0;
    1389: T504 = 1'h0;
    1390: T504 = 1'h0;
    1391: T504 = 1'h0;
    1392: T504 = 1'h0;
    1393: T504 = 1'h0;
    1394: T504 = 1'h0;
    1395: T504 = 1'h0;
    1396: T504 = 1'h0;
    1397: T504 = 1'h0;
    1398: T504 = 1'h0;
    1399: T504 = 1'h0;
    1400: T504 = 1'h0;
    1401: T504 = 1'h0;
    1402: T504 = 1'h0;
    1403: T504 = 1'h0;
    1404: T504 = 1'h0;
    1405: T504 = 1'h0;
    1406: T504 = 1'h0;
    1407: T504 = 1'h0;
    1408: T504 = 1'h0;
    1409: T504 = 1'h0;
    1410: T504 = 1'h0;
    1411: T504 = 1'h0;
    1412: T504 = 1'h0;
    1413: T504 = 1'h0;
    1414: T504 = 1'h0;
    1415: T504 = 1'h0;
    1416: T504 = 1'h0;
    1417: T504 = 1'h0;
    1418: T504 = 1'h0;
    1419: T504 = 1'h0;
    1420: T504 = 1'h0;
    1421: T504 = 1'h0;
    1422: T504 = 1'h0;
    1423: T504 = 1'h0;
    1424: T504 = 1'h0;
    1425: T504 = 1'h0;
    1426: T504 = 1'h0;
    1427: T504 = 1'h0;
    1428: T504 = 1'h0;
    1429: T504 = 1'h0;
    1430: T504 = 1'h0;
    1431: T504 = 1'h0;
    1432: T504 = 1'h0;
    1433: T504 = 1'h0;
    1434: T504 = 1'h0;
    1435: T504 = 1'h0;
    1436: T504 = 1'h0;
    1437: T504 = 1'h0;
    1438: T504 = 1'h0;
    1439: T504 = 1'h0;
    1440: T504 = 1'h0;
    1441: T504 = 1'h0;
    1442: T504 = 1'h0;
    1443: T504 = 1'h0;
    1444: T504 = 1'h0;
    1445: T504 = 1'h0;
    1446: T504 = 1'h0;
    1447: T504 = 1'h0;
    1448: T504 = 1'h0;
    1449: T504 = 1'h0;
    1450: T504 = 1'h0;
    1451: T504 = 1'h0;
    1452: T504 = 1'h0;
    1453: T504 = 1'h0;
    1454: T504 = 1'h0;
    1455: T504 = 1'h0;
    1456: T504 = 1'h0;
    1457: T504 = 1'h0;
    1458: T504 = 1'h0;
    1459: T504 = 1'h0;
    1460: T504 = 1'h0;
    1461: T504 = 1'h0;
    1462: T504 = 1'h0;
    1463: T504 = 1'h0;
    1464: T504 = 1'h0;
    1465: T504 = 1'h0;
    1466: T504 = 1'h0;
    1467: T504 = 1'h0;
    1468: T504 = 1'h0;
    1469: T504 = 1'h0;
    1470: T504 = 1'h0;
    1471: T504 = 1'h0;
    1472: T504 = 1'h0;
    1473: T504 = 1'h0;
    1474: T504 = 1'h0;
    1475: T504 = 1'h0;
    1476: T504 = 1'h0;
    1477: T504 = 1'h0;
    1478: T504 = 1'h0;
    1479: T504 = 1'h0;
    1480: T504 = 1'h0;
    1481: T504 = 1'h0;
    1482: T504 = 1'h0;
    1483: T504 = 1'h0;
    1484: T504 = 1'h0;
    1485: T504 = 1'h0;
    1486: T504 = 1'h0;
    1487: T504 = 1'h0;
    1488: T504 = 1'h0;
    1489: T504 = 1'h0;
    1490: T504 = 1'h0;
    1491: T504 = 1'h0;
    1492: T504 = 1'h0;
    1493: T504 = 1'h0;
    1494: T504 = 1'h0;
    1495: T504 = 1'h0;
    1496: T504 = 1'h0;
    1497: T504 = 1'h0;
    1498: T504 = 1'h0;
    1499: T504 = 1'h0;
    1500: T504 = 1'h0;
    1501: T504 = 1'h0;
    1502: T504 = 1'h0;
    1503: T504 = 1'h0;
    1504: T504 = 1'h0;
    1505: T504 = 1'h0;
    1506: T504 = 1'h0;
    1507: T504 = 1'h0;
    1508: T504 = 1'h0;
    1509: T504 = 1'h0;
    1510: T504 = 1'h0;
    1511: T504 = 1'h0;
    1512: T504 = 1'h0;
    1513: T504 = 1'h0;
    1514: T504 = 1'h0;
    1515: T504 = 1'h0;
    1516: T504 = 1'h0;
    1517: T504 = 1'h0;
    1518: T504 = 1'h0;
    1519: T504 = 1'h0;
    1520: T504 = 1'h0;
    1521: T504 = 1'h0;
    1522: T504 = 1'h0;
    1523: T504 = 1'h0;
    1524: T504 = 1'h0;
    1525: T504 = 1'h0;
    1526: T504 = 1'h0;
    1527: T504 = 1'h0;
    1528: T504 = 1'h0;
    1529: T504 = 1'h0;
    1530: T504 = 1'h0;
    1531: T504 = 1'h0;
    1532: T504 = 1'h0;
    1533: T504 = 1'h0;
    1534: T504 = 1'h0;
    1535: T504 = 1'h0;
    1536: T504 = 1'h0;
    1537: T504 = 1'h0;
    1538: T504 = 1'h0;
    1539: T504 = 1'h0;
    1540: T504 = 1'h0;
    1541: T504 = 1'h0;
    1542: T504 = 1'h0;
    1543: T504 = 1'h0;
    1544: T504 = 1'h0;
    1545: T504 = 1'h0;
    1546: T504 = 1'h0;
    1547: T504 = 1'h0;
    1548: T504 = 1'h0;
    1549: T504 = 1'h0;
    1550: T504 = 1'h0;
    1551: T504 = 1'h0;
    1552: T504 = 1'h0;
    1553: T504 = 1'h0;
    1554: T504 = 1'h0;
    1555: T504 = 1'h0;
    1556: T504 = 1'h0;
    1557: T504 = 1'h0;
    1558: T504 = 1'h0;
    1559: T504 = 1'h0;
    1560: T504 = 1'h0;
    1561: T504 = 1'h0;
    1562: T504 = 1'h0;
    1563: T504 = 1'h0;
    1564: T504 = 1'h0;
    1565: T504 = 1'h0;
    1566: T504 = 1'h0;
    1567: T504 = 1'h0;
    1568: T504 = 1'h0;
    1569: T504 = 1'h0;
    1570: T504 = 1'h0;
    1571: T504 = 1'h0;
    1572: T504 = 1'h0;
    1573: T504 = 1'h0;
    1574: T504 = 1'h0;
    1575: T504 = 1'h0;
    1576: T504 = 1'h0;
    1577: T504 = 1'h0;
    1578: T504 = 1'h0;
    1579: T504 = 1'h0;
    1580: T504 = 1'h0;
    1581: T504 = 1'h0;
    1582: T504 = 1'h0;
    1583: T504 = 1'h0;
    1584: T504 = 1'h0;
    1585: T504 = 1'h0;
    1586: T504 = 1'h0;
    1587: T504 = 1'h0;
    1588: T504 = 1'h0;
    1589: T504 = 1'h0;
    1590: T504 = 1'h0;
    1591: T504 = 1'h0;
    1592: T504 = 1'h0;
    1593: T504 = 1'h0;
    1594: T504 = 1'h0;
    1595: T504 = 1'h0;
    1596: T504 = 1'h0;
    1597: T504 = 1'h0;
    1598: T504 = 1'h0;
    1599: T504 = 1'h0;
    1600: T504 = 1'h0;
    1601: T504 = 1'h0;
    1602: T504 = 1'h0;
    1603: T504 = 1'h0;
    1604: T504 = 1'h0;
    1605: T504 = 1'h0;
    1606: T504 = 1'h0;
    1607: T504 = 1'h0;
    1608: T504 = 1'h0;
    1609: T504 = 1'h0;
    1610: T504 = 1'h0;
    1611: T504 = 1'h0;
    1612: T504 = 1'h0;
    1613: T504 = 1'h0;
    1614: T504 = 1'h0;
    1615: T504 = 1'h0;
    1616: T504 = 1'h0;
    1617: T504 = 1'h0;
    1618: T504 = 1'h0;
    1619: T504 = 1'h0;
    1620: T504 = 1'h0;
    1621: T504 = 1'h0;
    1622: T504 = 1'h0;
    1623: T504 = 1'h0;
    1624: T504 = 1'h0;
    1625: T504 = 1'h0;
    1626: T504 = 1'h0;
    1627: T504 = 1'h0;
    1628: T504 = 1'h0;
    1629: T504 = 1'h0;
    1630: T504 = 1'h0;
    1631: T504 = 1'h0;
    1632: T504 = 1'h0;
    1633: T504 = 1'h0;
    1634: T504 = 1'h0;
    1635: T504 = 1'h0;
    1636: T504 = 1'h0;
    1637: T504 = 1'h0;
    1638: T504 = 1'h0;
    1639: T504 = 1'h0;
    1640: T504 = 1'h0;
    1641: T504 = 1'h0;
    1642: T504 = 1'h0;
    1643: T504 = 1'h0;
    1644: T504 = 1'h0;
    1645: T504 = 1'h0;
    1646: T504 = 1'h0;
    1647: T504 = 1'h0;
    1648: T504 = 1'h0;
    1649: T504 = 1'h0;
    1650: T504 = 1'h0;
    1651: T504 = 1'h0;
    1652: T504 = 1'h0;
    1653: T504 = 1'h0;
    1654: T504 = 1'h0;
    1655: T504 = 1'h0;
    1656: T504 = 1'h0;
    1657: T504 = 1'h0;
    1658: T504 = 1'h0;
    1659: T504 = 1'h0;
    1660: T504 = 1'h0;
    1661: T504 = 1'h0;
    1662: T504 = 1'h0;
    1663: T504 = 1'h0;
    1664: T504 = 1'h0;
    1665: T504 = 1'h0;
    1666: T504 = 1'h0;
    1667: T504 = 1'h0;
    1668: T504 = 1'h0;
    1669: T504 = 1'h0;
    1670: T504 = 1'h0;
    1671: T504 = 1'h0;
    1672: T504 = 1'h0;
    1673: T504 = 1'h0;
    1674: T504 = 1'h0;
    1675: T504 = 1'h0;
    1676: T504 = 1'h0;
    1677: T504 = 1'h0;
    1678: T504 = 1'h0;
    1679: T504 = 1'h0;
    1680: T504 = 1'h0;
    1681: T504 = 1'h0;
    1682: T504 = 1'h0;
    1683: T504 = 1'h0;
    1684: T504 = 1'h0;
    1685: T504 = 1'h0;
    1686: T504 = 1'h0;
    1687: T504 = 1'h0;
    1688: T504 = 1'h0;
    1689: T504 = 1'h0;
    1690: T504 = 1'h0;
    1691: T504 = 1'h0;
    1692: T504 = 1'h0;
    1693: T504 = 1'h0;
    1694: T504 = 1'h0;
    1695: T504 = 1'h0;
    1696: T504 = 1'h0;
    1697: T504 = 1'h0;
    1698: T504 = 1'h0;
    1699: T504 = 1'h0;
    1700: T504 = 1'h0;
    1701: T504 = 1'h0;
    1702: T504 = 1'h0;
    1703: T504 = 1'h0;
    1704: T504 = 1'h0;
    1705: T504 = 1'h0;
    1706: T504 = 1'h0;
    1707: T504 = 1'h0;
    1708: T504 = 1'h0;
    1709: T504 = 1'h0;
    1710: T504 = 1'h0;
    1711: T504 = 1'h0;
    1712: T504 = 1'h0;
    1713: T504 = 1'h0;
    1714: T504 = 1'h0;
    1715: T504 = 1'h0;
    1716: T504 = 1'h0;
    1717: T504 = 1'h0;
    1718: T504 = 1'h0;
    1719: T504 = 1'h0;
    1720: T504 = 1'h0;
    1721: T504 = 1'h0;
    1722: T504 = 1'h0;
    1723: T504 = 1'h0;
    1724: T504 = 1'h0;
    1725: T504 = 1'h0;
    1726: T504 = 1'h0;
    1727: T504 = 1'h0;
    1728: T504 = 1'h0;
    1729: T504 = 1'h0;
    1730: T504 = 1'h0;
    1731: T504 = 1'h0;
    1732: T504 = 1'h0;
    1733: T504 = 1'h0;
    1734: T504 = 1'h0;
    1735: T504 = 1'h0;
    1736: T504 = 1'h0;
    1737: T504 = 1'h0;
    1738: T504 = 1'h0;
    1739: T504 = 1'h0;
    1740: T504 = 1'h0;
    1741: T504 = 1'h0;
    1742: T504 = 1'h0;
    1743: T504 = 1'h0;
    1744: T504 = 1'h0;
    1745: T504 = 1'h0;
    1746: T504 = 1'h0;
    1747: T504 = 1'h0;
    1748: T504 = 1'h0;
    1749: T504 = 1'h0;
    1750: T504 = 1'h0;
    1751: T504 = 1'h0;
    1752: T504 = 1'h0;
    1753: T504 = 1'h0;
    1754: T504 = 1'h0;
    1755: T504 = 1'h0;
    1756: T504 = 1'h0;
    1757: T504 = 1'h0;
    1758: T504 = 1'h0;
    1759: T504 = 1'h0;
    1760: T504 = 1'h0;
    1761: T504 = 1'h0;
    1762: T504 = 1'h0;
    1763: T504 = 1'h0;
    1764: T504 = 1'h0;
    1765: T504 = 1'h0;
    1766: T504 = 1'h0;
    1767: T504 = 1'h0;
    1768: T504 = 1'h0;
    1769: T504 = 1'h0;
    1770: T504 = 1'h0;
    1771: T504 = 1'h0;
    1772: T504 = 1'h0;
    1773: T504 = 1'h0;
    1774: T504 = 1'h0;
    1775: T504 = 1'h0;
    1776: T504 = 1'h0;
    1777: T504 = 1'h0;
    1778: T504 = 1'h0;
    1779: T504 = 1'h0;
    1780: T504 = 1'h0;
    1781: T504 = 1'h0;
    1782: T504 = 1'h0;
    1783: T504 = 1'h0;
    1784: T504 = 1'h0;
    1785: T504 = 1'h0;
    1786: T504 = 1'h0;
    1787: T504 = 1'h0;
    1788: T504 = 1'h0;
    1789: T504 = 1'h0;
    1790: T504 = 1'h0;
    1791: T504 = 1'h0;
    1792: T504 = 1'h0;
    1793: T504 = 1'h0;
    1794: T504 = 1'h0;
    1795: T504 = 1'h0;
    1796: T504 = 1'h0;
    1797: T504 = 1'h0;
    1798: T504 = 1'h0;
    1799: T504 = 1'h0;
    1800: T504 = 1'h0;
    1801: T504 = 1'h0;
    1802: T504 = 1'h0;
    1803: T504 = 1'h0;
    1804: T504 = 1'h0;
    1805: T504 = 1'h0;
    1806: T504 = 1'h0;
    1807: T504 = 1'h0;
    1808: T504 = 1'h0;
    1809: T504 = 1'h0;
    1810: T504 = 1'h0;
    1811: T504 = 1'h0;
    1812: T504 = 1'h0;
    1813: T504 = 1'h0;
    1814: T504 = 1'h0;
    1815: T504 = 1'h0;
    1816: T504 = 1'h0;
    1817: T504 = 1'h0;
    1818: T504 = 1'h0;
    1819: T504 = 1'h0;
    1820: T504 = 1'h0;
    1821: T504 = 1'h0;
    1822: T504 = 1'h0;
    1823: T504 = 1'h0;
    1824: T504 = 1'h0;
    1825: T504 = 1'h0;
    1826: T504 = 1'h0;
    1827: T504 = 1'h0;
    1828: T504 = 1'h0;
    1829: T504 = 1'h0;
    1830: T504 = 1'h0;
    1831: T504 = 1'h0;
    1832: T504 = 1'h0;
    1833: T504 = 1'h0;
    1834: T504 = 1'h0;
    1835: T504 = 1'h0;
    1836: T504 = 1'h0;
    1837: T504 = 1'h0;
    1838: T504 = 1'h0;
    1839: T504 = 1'h0;
    1840: T504 = 1'h0;
    1841: T504 = 1'h0;
    1842: T504 = 1'h0;
    1843: T504 = 1'h0;
    1844: T504 = 1'h0;
    1845: T504 = 1'h0;
    1846: T504 = 1'h0;
    1847: T504 = 1'h0;
    1848: T504 = 1'h0;
    1849: T504 = 1'h0;
    1850: T504 = 1'h0;
    1851: T504 = 1'h0;
    1852: T504 = 1'h0;
    1853: T504 = 1'h0;
    1854: T504 = 1'h0;
    1855: T504 = 1'h0;
    1856: T504 = 1'h0;
    1857: T504 = 1'h0;
    1858: T504 = 1'h0;
    1859: T504 = 1'h0;
    1860: T504 = 1'h0;
    1861: T504 = 1'h0;
    1862: T504 = 1'h0;
    1863: T504 = 1'h0;
    1864: T504 = 1'h0;
    1865: T504 = 1'h0;
    1866: T504 = 1'h0;
    1867: T504 = 1'h0;
    1868: T504 = 1'h0;
    1869: T504 = 1'h0;
    1870: T504 = 1'h0;
    1871: T504 = 1'h0;
    1872: T504 = 1'h0;
    1873: T504 = 1'h0;
    1874: T504 = 1'h0;
    1875: T504 = 1'h0;
    1876: T504 = 1'h0;
    1877: T504 = 1'h0;
    1878: T504 = 1'h0;
    1879: T504 = 1'h0;
    1880: T504 = 1'h0;
    1881: T504 = 1'h0;
    1882: T504 = 1'h0;
    1883: T504 = 1'h0;
    1884: T504 = 1'h0;
    1885: T504 = 1'h0;
    1886: T504 = 1'h0;
    1887: T504 = 1'h0;
    1888: T504 = 1'h0;
    1889: T504 = 1'h0;
    1890: T504 = 1'h0;
    1891: T504 = 1'h0;
    1892: T504 = 1'h0;
    1893: T504 = 1'h0;
    1894: T504 = 1'h0;
    1895: T504 = 1'h0;
    1896: T504 = 1'h0;
    1897: T504 = 1'h0;
    1898: T504 = 1'h0;
    1899: T504 = 1'h0;
    1900: T504 = 1'h0;
    1901: T504 = 1'h0;
    1902: T504 = 1'h0;
    1903: T504 = 1'h0;
    1904: T504 = 1'h0;
    1905: T504 = 1'h0;
    1906: T504 = 1'h0;
    1907: T504 = 1'h0;
    1908: T504 = 1'h0;
    1909: T504 = 1'h0;
    1910: T504 = 1'h0;
    1911: T504 = 1'h0;
    1912: T504 = 1'h0;
    1913: T504 = 1'h0;
    1914: T504 = 1'h0;
    1915: T504 = 1'h0;
    1916: T504 = 1'h0;
    1917: T504 = 1'h0;
    1918: T504 = 1'h0;
    1919: T504 = 1'h0;
    1920: T504 = 1'h0;
    1921: T504 = 1'h0;
    1922: T504 = 1'h0;
    1923: T504 = 1'h0;
    1924: T504 = 1'h0;
    1925: T504 = 1'h0;
    1926: T504 = 1'h0;
    1927: T504 = 1'h0;
    1928: T504 = 1'h0;
    1929: T504 = 1'h0;
    1930: T504 = 1'h0;
    1931: T504 = 1'h0;
    1932: T504 = 1'h0;
    1933: T504 = 1'h0;
    1934: T504 = 1'h0;
    1935: T504 = 1'h0;
    1936: T504 = 1'h0;
    1937: T504 = 1'h0;
    1938: T504 = 1'h0;
    1939: T504 = 1'h0;
    1940: T504 = 1'h0;
    1941: T504 = 1'h0;
    1942: T504 = 1'h0;
    1943: T504 = 1'h0;
    1944: T504 = 1'h0;
    1945: T504 = 1'h0;
    1946: T504 = 1'h0;
    1947: T504 = 1'h0;
    1948: T504 = 1'h0;
    1949: T504 = 1'h0;
    1950: T504 = 1'h0;
    1951: T504 = 1'h0;
    1952: T504 = 1'h0;
    1953: T504 = 1'h0;
    1954: T504 = 1'h0;
    1955: T504 = 1'h0;
    1956: T504 = 1'h0;
    1957: T504 = 1'h0;
    1958: T504 = 1'h0;
    1959: T504 = 1'h0;
    1960: T504 = 1'h0;
    1961: T504 = 1'h0;
    1962: T504 = 1'h0;
    1963: T504 = 1'h0;
    1964: T504 = 1'h0;
    1965: T504 = 1'h0;
    1966: T504 = 1'h0;
    1967: T504 = 1'h0;
    1968: T504 = 1'h0;
    1969: T504 = 1'h0;
    1970: T504 = 1'h0;
    1971: T504 = 1'h0;
    1972: T504 = 1'h0;
    1973: T504 = 1'h0;
    1974: T504 = 1'h0;
    1975: T504 = 1'h0;
    1976: T504 = 1'h0;
    1977: T504 = 1'h0;
    1978: T504 = 1'h0;
    1979: T504 = 1'h0;
    1980: T504 = 1'h0;
    1981: T504 = 1'h0;
    1982: T504 = 1'h0;
    1983: T504 = 1'h0;
    1984: T504 = 1'h0;
    1985: T504 = 1'h0;
    1986: T504 = 1'h0;
    1987: T504 = 1'h0;
    1988: T504 = 1'h0;
    1989: T504 = 1'h0;
    1990: T504 = 1'h0;
    1991: T504 = 1'h0;
    1992: T504 = 1'h0;
    1993: T504 = 1'h0;
    1994: T504 = 1'h0;
    1995: T504 = 1'h0;
    1996: T504 = 1'h0;
    1997: T504 = 1'h0;
    1998: T504 = 1'h0;
    1999: T504 = 1'h0;
    2000: T504 = 1'h0;
    2001: T504 = 1'h0;
    2002: T504 = 1'h0;
    2003: T504 = 1'h0;
    2004: T504 = 1'h0;
    2005: T504 = 1'h0;
    2006: T504 = 1'h0;
    2007: T504 = 1'h0;
    2008: T504 = 1'h0;
    2009: T504 = 1'h0;
    2010: T504 = 1'h0;
    2011: T504 = 1'h0;
    2012: T504 = 1'h0;
    2013: T504 = 1'h0;
    2014: T504 = 1'h0;
    2015: T504 = 1'h0;
    2016: T504 = 1'h0;
    2017: T504 = 1'h0;
    2018: T504 = 1'h0;
    2019: T504 = 1'h0;
    2020: T504 = 1'h0;
    2021: T504 = 1'h0;
    2022: T504 = 1'h0;
    2023: T504 = 1'h0;
    2024: T504 = 1'h0;
    2025: T504 = 1'h0;
    2026: T504 = 1'h0;
    2027: T504 = 1'h0;
    2028: T504 = 1'h0;
    2029: T504 = 1'h0;
    2030: T504 = 1'h0;
    2031: T504 = 1'h0;
    2032: T504 = 1'h0;
    2033: T504 = 1'h0;
    2034: T504 = 1'h0;
    2035: T504 = 1'h0;
    2036: T504 = 1'h0;
    2037: T504 = 1'h0;
    2038: T504 = 1'h0;
    2039: T504 = 1'h0;
    2040: T504 = 1'h0;
    2041: T504 = 1'h0;
    2042: T504 = 1'h0;
    2043: T504 = 1'h0;
    2044: T504 = 1'h0;
    2045: T504 = 1'h0;
    2046: T504 = 1'h0;
    2047: T504 = 1'h0;
    2048: T504 = 1'h0;
    2049: T504 = 1'h0;
    2050: T504 = 1'h0;
    2051: T504 = 1'h0;
    2052: T504 = 1'h0;
    2053: T504 = 1'h0;
    2054: T504 = 1'h0;
    2055: T504 = 1'h0;
    2056: T504 = 1'h0;
    2057: T504 = 1'h0;
    2058: T504 = 1'h0;
    2059: T504 = 1'h0;
    2060: T504 = 1'h0;
    2061: T504 = 1'h0;
    2062: T504 = 1'h0;
    2063: T504 = 1'h0;
    2064: T504 = 1'h0;
    2065: T504 = 1'h0;
    2066: T504 = 1'h0;
    2067: T504 = 1'h0;
    2068: T504 = 1'h0;
    2069: T504 = 1'h0;
    2070: T504 = 1'h0;
    2071: T504 = 1'h0;
    2072: T504 = 1'h0;
    2073: T504 = 1'h0;
    2074: T504 = 1'h0;
    2075: T504 = 1'h0;
    2076: T504 = 1'h0;
    2077: T504 = 1'h0;
    2078: T504 = 1'h0;
    2079: T504 = 1'h0;
    2080: T504 = 1'h0;
    2081: T504 = 1'h0;
    2082: T504 = 1'h0;
    2083: T504 = 1'h0;
    2084: T504 = 1'h0;
    2085: T504 = 1'h0;
    2086: T504 = 1'h0;
    2087: T504 = 1'h0;
    2088: T504 = 1'h0;
    2089: T504 = 1'h0;
    2090: T504 = 1'h0;
    2091: T504 = 1'h0;
    2092: T504 = 1'h0;
    2093: T504 = 1'h0;
    2094: T504 = 1'h0;
    2095: T504 = 1'h0;
    2096: T504 = 1'h0;
    2097: T504 = 1'h0;
    2098: T504 = 1'h0;
    2099: T504 = 1'h0;
    2100: T504 = 1'h0;
    2101: T504 = 1'h0;
    2102: T504 = 1'h0;
    2103: T504 = 1'h0;
    2104: T504 = 1'h0;
    2105: T504 = 1'h0;
    2106: T504 = 1'h0;
    2107: T504 = 1'h0;
    2108: T504 = 1'h0;
    2109: T504 = 1'h0;
    2110: T504 = 1'h0;
    2111: T504 = 1'h0;
    2112: T504 = 1'h0;
    2113: T504 = 1'h0;
    2114: T504 = 1'h0;
    2115: T504 = 1'h0;
    2116: T504 = 1'h0;
    2117: T504 = 1'h0;
    2118: T504 = 1'h0;
    2119: T504 = 1'h0;
    2120: T504 = 1'h0;
    2121: T504 = 1'h0;
    2122: T504 = 1'h0;
    2123: T504 = 1'h0;
    2124: T504 = 1'h0;
    2125: T504 = 1'h0;
    2126: T504 = 1'h0;
    2127: T504 = 1'h0;
    2128: T504 = 1'h0;
    2129: T504 = 1'h0;
    2130: T504 = 1'h0;
    2131: T504 = 1'h0;
    2132: T504 = 1'h0;
    2133: T504 = 1'h0;
    2134: T504 = 1'h0;
    2135: T504 = 1'h0;
    2136: T504 = 1'h0;
    2137: T504 = 1'h0;
    2138: T504 = 1'h0;
    2139: T504 = 1'h0;
    2140: T504 = 1'h0;
    2141: T504 = 1'h0;
    2142: T504 = 1'h0;
    2143: T504 = 1'h0;
    2144: T504 = 1'h0;
    2145: T504 = 1'h0;
    2146: T504 = 1'h0;
    2147: T504 = 1'h0;
    2148: T504 = 1'h0;
    2149: T504 = 1'h0;
    2150: T504 = 1'h0;
    2151: T504 = 1'h0;
    2152: T504 = 1'h0;
    2153: T504 = 1'h0;
    2154: T504 = 1'h0;
    2155: T504 = 1'h0;
    2156: T504 = 1'h0;
    2157: T504 = 1'h0;
    2158: T504 = 1'h0;
    2159: T504 = 1'h0;
    2160: T504 = 1'h0;
    2161: T504 = 1'h0;
    2162: T504 = 1'h0;
    2163: T504 = 1'h0;
    2164: T504 = 1'h0;
    2165: T504 = 1'h0;
    2166: T504 = 1'h0;
    2167: T504 = 1'h0;
    2168: T504 = 1'h0;
    2169: T504 = 1'h0;
    2170: T504 = 1'h0;
    2171: T504 = 1'h0;
    2172: T504 = 1'h0;
    2173: T504 = 1'h0;
    2174: T504 = 1'h0;
    2175: T504 = 1'h0;
    2176: T504 = 1'h0;
    2177: T504 = 1'h0;
    2178: T504 = 1'h0;
    2179: T504 = 1'h0;
    2180: T504 = 1'h0;
    2181: T504 = 1'h0;
    2182: T504 = 1'h0;
    2183: T504 = 1'h0;
    2184: T504 = 1'h0;
    2185: T504 = 1'h0;
    2186: T504 = 1'h0;
    2187: T504 = 1'h0;
    2188: T504 = 1'h0;
    2189: T504 = 1'h0;
    2190: T504 = 1'h0;
    2191: T504 = 1'h0;
    2192: T504 = 1'h0;
    2193: T504 = 1'h0;
    2194: T504 = 1'h0;
    2195: T504 = 1'h0;
    2196: T504 = 1'h0;
    2197: T504 = 1'h0;
    2198: T504 = 1'h0;
    2199: T504 = 1'h0;
    2200: T504 = 1'h0;
    2201: T504 = 1'h0;
    2202: T504 = 1'h0;
    2203: T504 = 1'h0;
    2204: T504 = 1'h0;
    2205: T504 = 1'h0;
    2206: T504 = 1'h0;
    2207: T504 = 1'h0;
    2208: T504 = 1'h0;
    2209: T504 = 1'h0;
    2210: T504 = 1'h0;
    2211: T504 = 1'h0;
    2212: T504 = 1'h0;
    2213: T504 = 1'h0;
    2214: T504 = 1'h0;
    2215: T504 = 1'h0;
    2216: T504 = 1'h0;
    2217: T504 = 1'h0;
    2218: T504 = 1'h0;
    2219: T504 = 1'h0;
    2220: T504 = 1'h0;
    2221: T504 = 1'h0;
    2222: T504 = 1'h0;
    2223: T504 = 1'h0;
    2224: T504 = 1'h0;
    2225: T504 = 1'h0;
    2226: T504 = 1'h0;
    2227: T504 = 1'h0;
    2228: T504 = 1'h0;
    2229: T504 = 1'h0;
    2230: T504 = 1'h0;
    2231: T504 = 1'h0;
    2232: T504 = 1'h0;
    2233: T504 = 1'h0;
    2234: T504 = 1'h0;
    2235: T504 = 1'h0;
    2236: T504 = 1'h0;
    2237: T504 = 1'h0;
    2238: T504 = 1'h0;
    2239: T504 = 1'h0;
    2240: T504 = 1'h0;
    2241: T504 = 1'h0;
    2242: T504 = 1'h0;
    2243: T504 = 1'h0;
    2244: T504 = 1'h0;
    2245: T504 = 1'h0;
    2246: T504 = 1'h0;
    2247: T504 = 1'h0;
    2248: T504 = 1'h0;
    2249: T504 = 1'h0;
    2250: T504 = 1'h0;
    2251: T504 = 1'h0;
    2252: T504 = 1'h0;
    2253: T504 = 1'h0;
    2254: T504 = 1'h0;
    2255: T504 = 1'h0;
    2256: T504 = 1'h0;
    2257: T504 = 1'h0;
    2258: T504 = 1'h0;
    2259: T504 = 1'h0;
    2260: T504 = 1'h0;
    2261: T504 = 1'h0;
    2262: T504 = 1'h0;
    2263: T504 = 1'h0;
    2264: T504 = 1'h0;
    2265: T504 = 1'h0;
    2266: T504 = 1'h0;
    2267: T504 = 1'h0;
    2268: T504 = 1'h0;
    2269: T504 = 1'h0;
    2270: T504 = 1'h0;
    2271: T504 = 1'h0;
    2272: T504 = 1'h0;
    2273: T504 = 1'h0;
    2274: T504 = 1'h0;
    2275: T504 = 1'h0;
    2276: T504 = 1'h0;
    2277: T504 = 1'h0;
    2278: T504 = 1'h0;
    2279: T504 = 1'h0;
    2280: T504 = 1'h0;
    2281: T504 = 1'h0;
    2282: T504 = 1'h0;
    2283: T504 = 1'h0;
    2284: T504 = 1'h0;
    2285: T504 = 1'h0;
    2286: T504 = 1'h0;
    2287: T504 = 1'h0;
    2288: T504 = 1'h0;
    2289: T504 = 1'h0;
    2290: T504 = 1'h0;
    2291: T504 = 1'h0;
    2292: T504 = 1'h0;
    2293: T504 = 1'h0;
    2294: T504 = 1'h0;
    2295: T504 = 1'h0;
    2296: T504 = 1'h0;
    2297: T504 = 1'h0;
    2298: T504 = 1'h0;
    2299: T504 = 1'h0;
    2300: T504 = 1'h0;
    2301: T504 = 1'h0;
    2302: T504 = 1'h0;
    2303: T504 = 1'h0;
    2304: T504 = 1'h0;
    2305: T504 = 1'h0;
    2306: T504 = 1'h0;
    2307: T504 = 1'h0;
    2308: T504 = 1'h0;
    2309: T504 = 1'h0;
    2310: T504 = 1'h0;
    2311: T504 = 1'h0;
    2312: T504 = 1'h0;
    2313: T504 = 1'h0;
    2314: T504 = 1'h0;
    2315: T504 = 1'h0;
    2316: T504 = 1'h0;
    2317: T504 = 1'h0;
    2318: T504 = 1'h0;
    2319: T504 = 1'h0;
    2320: T504 = 1'h0;
    2321: T504 = 1'h0;
    2322: T504 = 1'h0;
    2323: T504 = 1'h0;
    2324: T504 = 1'h0;
    2325: T504 = 1'h0;
    2326: T504 = 1'h0;
    2327: T504 = 1'h0;
    2328: T504 = 1'h0;
    2329: T504 = 1'h0;
    2330: T504 = 1'h0;
    2331: T504 = 1'h0;
    2332: T504 = 1'h0;
    2333: T504 = 1'h0;
    2334: T504 = 1'h0;
    2335: T504 = 1'h0;
    2336: T504 = 1'h0;
    2337: T504 = 1'h0;
    2338: T504 = 1'h0;
    2339: T504 = 1'h0;
    2340: T504 = 1'h0;
    2341: T504 = 1'h0;
    2342: T504 = 1'h0;
    2343: T504 = 1'h0;
    2344: T504 = 1'h0;
    2345: T504 = 1'h0;
    2346: T504 = 1'h0;
    2347: T504 = 1'h0;
    2348: T504 = 1'h0;
    2349: T504 = 1'h0;
    2350: T504 = 1'h0;
    2351: T504 = 1'h0;
    2352: T504 = 1'h0;
    2353: T504 = 1'h0;
    2354: T504 = 1'h0;
    2355: T504 = 1'h0;
    2356: T504 = 1'h0;
    2357: T504 = 1'h0;
    2358: T504 = 1'h0;
    2359: T504 = 1'h0;
    2360: T504 = 1'h0;
    2361: T504 = 1'h0;
    2362: T504 = 1'h0;
    2363: T504 = 1'h0;
    2364: T504 = 1'h0;
    2365: T504 = 1'h0;
    2366: T504 = 1'h0;
    2367: T504 = 1'h0;
    2368: T504 = 1'h0;
    2369: T504 = 1'h0;
    2370: T504 = 1'h0;
    2371: T504 = 1'h0;
    2372: T504 = 1'h0;
    2373: T504 = 1'h0;
    2374: T504 = 1'h0;
    2375: T504 = 1'h0;
    2376: T504 = 1'h0;
    2377: T504 = 1'h0;
    2378: T504 = 1'h0;
    2379: T504 = 1'h0;
    2380: T504 = 1'h0;
    2381: T504 = 1'h0;
    2382: T504 = 1'h0;
    2383: T504 = 1'h0;
    2384: T504 = 1'h0;
    2385: T504 = 1'h0;
    2386: T504 = 1'h0;
    2387: T504 = 1'h0;
    2388: T504 = 1'h0;
    2389: T504 = 1'h0;
    2390: T504 = 1'h0;
    2391: T504 = 1'h0;
    2392: T504 = 1'h0;
    2393: T504 = 1'h0;
    2394: T504 = 1'h0;
    2395: T504 = 1'h0;
    2396: T504 = 1'h0;
    2397: T504 = 1'h0;
    2398: T504 = 1'h0;
    2399: T504 = 1'h0;
    2400: T504 = 1'h0;
    2401: T504 = 1'h0;
    2402: T504 = 1'h0;
    2403: T504 = 1'h0;
    2404: T504 = 1'h0;
    2405: T504 = 1'h0;
    2406: T504 = 1'h0;
    2407: T504 = 1'h0;
    2408: T504 = 1'h0;
    2409: T504 = 1'h0;
    2410: T504 = 1'h0;
    2411: T504 = 1'h0;
    2412: T504 = 1'h0;
    2413: T504 = 1'h0;
    2414: T504 = 1'h0;
    2415: T504 = 1'h0;
    2416: T504 = 1'h0;
    2417: T504 = 1'h0;
    2418: T504 = 1'h0;
    2419: T504 = 1'h0;
    2420: T504 = 1'h0;
    2421: T504 = 1'h0;
    2422: T504 = 1'h0;
    2423: T504 = 1'h0;
    2424: T504 = 1'h0;
    2425: T504 = 1'h0;
    2426: T504 = 1'h0;
    2427: T504 = 1'h0;
    2428: T504 = 1'h0;
    2429: T504 = 1'h0;
    2430: T504 = 1'h0;
    2431: T504 = 1'h0;
    2432: T504 = 1'h0;
    2433: T504 = 1'h0;
    2434: T504 = 1'h0;
    2435: T504 = 1'h0;
    2436: T504 = 1'h0;
    2437: T504 = 1'h0;
    2438: T504 = 1'h0;
    2439: T504 = 1'h0;
    2440: T504 = 1'h0;
    2441: T504 = 1'h0;
    2442: T504 = 1'h0;
    2443: T504 = 1'h0;
    2444: T504 = 1'h0;
    2445: T504 = 1'h0;
    2446: T504 = 1'h0;
    2447: T504 = 1'h0;
    2448: T504 = 1'h0;
    2449: T504 = 1'h0;
    2450: T504 = 1'h0;
    2451: T504 = 1'h0;
    2452: T504 = 1'h0;
    2453: T504 = 1'h0;
    2454: T504 = 1'h0;
    2455: T504 = 1'h0;
    2456: T504 = 1'h0;
    2457: T504 = 1'h0;
    2458: T504 = 1'h0;
    2459: T504 = 1'h0;
    2460: T504 = 1'h0;
    2461: T504 = 1'h0;
    2462: T504 = 1'h0;
    2463: T504 = 1'h0;
    2464: T504 = 1'h0;
    2465: T504 = 1'h0;
    2466: T504 = 1'h0;
    2467: T504 = 1'h0;
    2468: T504 = 1'h0;
    2469: T504 = 1'h0;
    2470: T504 = 1'h0;
    2471: T504 = 1'h0;
    2472: T504 = 1'h0;
    2473: T504 = 1'h0;
    2474: T504 = 1'h0;
    2475: T504 = 1'h0;
    2476: T504 = 1'h0;
    2477: T504 = 1'h0;
    2478: T504 = 1'h0;
    2479: T504 = 1'h0;
    2480: T504 = 1'h0;
    2481: T504 = 1'h0;
    2482: T504 = 1'h0;
    2483: T504 = 1'h0;
    2484: T504 = 1'h0;
    2485: T504 = 1'h0;
    2486: T504 = 1'h0;
    2487: T504 = 1'h0;
    2488: T504 = 1'h0;
    2489: T504 = 1'h0;
    2490: T504 = 1'h0;
    2491: T504 = 1'h0;
    2492: T504 = 1'h0;
    2493: T504 = 1'h0;
    2494: T504 = 1'h0;
    2495: T504 = 1'h0;
    2496: T504 = 1'h0;
    2497: T504 = 1'h0;
    2498: T504 = 1'h0;
    2499: T504 = 1'h0;
    2500: T504 = 1'h0;
    2501: T504 = 1'h0;
    2502: T504 = 1'h0;
    2503: T504 = 1'h0;
    2504: T504 = 1'h0;
    2505: T504 = 1'h0;
    2506: T504 = 1'h0;
    2507: T504 = 1'h0;
    2508: T504 = 1'h0;
    2509: T504 = 1'h0;
    2510: T504 = 1'h0;
    2511: T504 = 1'h0;
    2512: T504 = 1'h0;
    2513: T504 = 1'h0;
    2514: T504 = 1'h0;
    2515: T504 = 1'h0;
    2516: T504 = 1'h0;
    2517: T504 = 1'h0;
    2518: T504 = 1'h0;
    2519: T504 = 1'h0;
    2520: T504 = 1'h0;
    2521: T504 = 1'h0;
    2522: T504 = 1'h0;
    2523: T504 = 1'h0;
    2524: T504 = 1'h0;
    2525: T504 = 1'h0;
    2526: T504 = 1'h0;
    2527: T504 = 1'h0;
    2528: T504 = 1'h0;
    2529: T504 = 1'h0;
    2530: T504 = 1'h0;
    2531: T504 = 1'h0;
    2532: T504 = 1'h0;
    2533: T504 = 1'h0;
    2534: T504 = 1'h0;
    2535: T504 = 1'h0;
    2536: T504 = 1'h0;
    2537: T504 = 1'h0;
    2538: T504 = 1'h0;
    2539: T504 = 1'h0;
    2540: T504 = 1'h0;
    2541: T504 = 1'h0;
    2542: T504 = 1'h0;
    2543: T504 = 1'h0;
    2544: T504 = 1'h0;
    2545: T504 = 1'h0;
    2546: T504 = 1'h0;
    2547: T504 = 1'h0;
    2548: T504 = 1'h0;
    2549: T504 = 1'h0;
    2550: T504 = 1'h0;
    2551: T504 = 1'h0;
    2552: T504 = 1'h0;
    2553: T504 = 1'h0;
    2554: T504 = 1'h0;
    2555: T504 = 1'h0;
    2556: T504 = 1'h0;
    2557: T504 = 1'h0;
    2558: T504 = 1'h0;
    2559: T504 = 1'h0;
    2560: T504 = 1'h0;
    2561: T504 = 1'h0;
    2562: T504 = 1'h0;
    2563: T504 = 1'h0;
    2564: T504 = 1'h0;
    2565: T504 = 1'h0;
    2566: T504 = 1'h0;
    2567: T504 = 1'h0;
    2568: T504 = 1'h0;
    2569: T504 = 1'h0;
    2570: T504 = 1'h0;
    2571: T504 = 1'h0;
    2572: T504 = 1'h0;
    2573: T504 = 1'h0;
    2574: T504 = 1'h0;
    2575: T504 = 1'h0;
    2576: T504 = 1'h0;
    2577: T504 = 1'h0;
    2578: T504 = 1'h0;
    2579: T504 = 1'h0;
    2580: T504 = 1'h0;
    2581: T504 = 1'h0;
    2582: T504 = 1'h0;
    2583: T504 = 1'h0;
    2584: T504 = 1'h0;
    2585: T504 = 1'h0;
    2586: T504 = 1'h0;
    2587: T504 = 1'h0;
    2588: T504 = 1'h0;
    2589: T504 = 1'h0;
    2590: T504 = 1'h0;
    2591: T504 = 1'h0;
    2592: T504 = 1'h0;
    2593: T504 = 1'h0;
    2594: T504 = 1'h0;
    2595: T504 = 1'h0;
    2596: T504 = 1'h0;
    2597: T504 = 1'h0;
    2598: T504 = 1'h0;
    2599: T504 = 1'h0;
    2600: T504 = 1'h0;
    2601: T504 = 1'h0;
    2602: T504 = 1'h0;
    2603: T504 = 1'h0;
    2604: T504 = 1'h0;
    2605: T504 = 1'h0;
    2606: T504 = 1'h0;
    2607: T504 = 1'h0;
    2608: T504 = 1'h0;
    2609: T504 = 1'h0;
    2610: T504 = 1'h0;
    2611: T504 = 1'h0;
    2612: T504 = 1'h0;
    2613: T504 = 1'h0;
    2614: T504 = 1'h0;
    2615: T504 = 1'h0;
    2616: T504 = 1'h0;
    2617: T504 = 1'h0;
    2618: T504 = 1'h0;
    2619: T504 = 1'h0;
    2620: T504 = 1'h0;
    2621: T504 = 1'h0;
    2622: T504 = 1'h0;
    2623: T504 = 1'h0;
    2624: T504 = 1'h0;
    2625: T504 = 1'h0;
    2626: T504 = 1'h0;
    2627: T504 = 1'h0;
    2628: T504 = 1'h0;
    2629: T504 = 1'h0;
    2630: T504 = 1'h0;
    2631: T504 = 1'h0;
    2632: T504 = 1'h0;
    2633: T504 = 1'h0;
    2634: T504 = 1'h0;
    2635: T504 = 1'h0;
    2636: T504 = 1'h0;
    2637: T504 = 1'h0;
    2638: T504 = 1'h0;
    2639: T504 = 1'h0;
    2640: T504 = 1'h0;
    2641: T504 = 1'h0;
    2642: T504 = 1'h0;
    2643: T504 = 1'h0;
    2644: T504 = 1'h0;
    2645: T504 = 1'h0;
    2646: T504 = 1'h0;
    2647: T504 = 1'h0;
    2648: T504 = 1'h0;
    2649: T504 = 1'h0;
    2650: T504 = 1'h0;
    2651: T504 = 1'h0;
    2652: T504 = 1'h0;
    2653: T504 = 1'h0;
    2654: T504 = 1'h0;
    2655: T504 = 1'h0;
    2656: T504 = 1'h0;
    2657: T504 = 1'h0;
    2658: T504 = 1'h0;
    2659: T504 = 1'h0;
    2660: T504 = 1'h0;
    2661: T504 = 1'h0;
    2662: T504 = 1'h0;
    2663: T504 = 1'h0;
    2664: T504 = 1'h0;
    2665: T504 = 1'h0;
    2666: T504 = 1'h0;
    2667: T504 = 1'h0;
    2668: T504 = 1'h0;
    2669: T504 = 1'h0;
    2670: T504 = 1'h0;
    2671: T504 = 1'h0;
    2672: T504 = 1'h0;
    2673: T504 = 1'h0;
    2674: T504 = 1'h0;
    2675: T504 = 1'h0;
    2676: T504 = 1'h0;
    2677: T504 = 1'h0;
    2678: T504 = 1'h0;
    2679: T504 = 1'h0;
    2680: T504 = 1'h0;
    2681: T504 = 1'h0;
    2682: T504 = 1'h0;
    2683: T504 = 1'h0;
    2684: T504 = 1'h0;
    2685: T504 = 1'h0;
    2686: T504 = 1'h0;
    2687: T504 = 1'h0;
    2688: T504 = 1'h0;
    2689: T504 = 1'h0;
    2690: T504 = 1'h0;
    2691: T504 = 1'h0;
    2692: T504 = 1'h0;
    2693: T504 = 1'h0;
    2694: T504 = 1'h0;
    2695: T504 = 1'h0;
    2696: T504 = 1'h0;
    2697: T504 = 1'h0;
    2698: T504 = 1'h0;
    2699: T504 = 1'h0;
    2700: T504 = 1'h0;
    2701: T504 = 1'h0;
    2702: T504 = 1'h0;
    2703: T504 = 1'h0;
    2704: T504 = 1'h0;
    2705: T504 = 1'h0;
    2706: T504 = 1'h0;
    2707: T504 = 1'h0;
    2708: T504 = 1'h0;
    2709: T504 = 1'h0;
    2710: T504 = 1'h0;
    2711: T504 = 1'h0;
    2712: T504 = 1'h0;
    2713: T504 = 1'h0;
    2714: T504 = 1'h0;
    2715: T504 = 1'h0;
    2716: T504 = 1'h0;
    2717: T504 = 1'h0;
    2718: T504 = 1'h0;
    2719: T504 = 1'h0;
    2720: T504 = 1'h0;
    2721: T504 = 1'h0;
    2722: T504 = 1'h0;
    2723: T504 = 1'h0;
    2724: T504 = 1'h0;
    2725: T504 = 1'h0;
    2726: T504 = 1'h0;
    2727: T504 = 1'h0;
    2728: T504 = 1'h0;
    2729: T504 = 1'h0;
    2730: T504 = 1'h0;
    2731: T504 = 1'h0;
    2732: T504 = 1'h0;
    2733: T504 = 1'h0;
    2734: T504 = 1'h0;
    2735: T504 = 1'h0;
    2736: T504 = 1'h0;
    2737: T504 = 1'h0;
    2738: T504 = 1'h0;
    2739: T504 = 1'h0;
    2740: T504 = 1'h0;
    2741: T504 = 1'h0;
    2742: T504 = 1'h0;
    2743: T504 = 1'h0;
    2744: T504 = 1'h0;
    2745: T504 = 1'h0;
    2746: T504 = 1'h0;
    2747: T504 = 1'h0;
    2748: T504 = 1'h0;
    2749: T504 = 1'h0;
    2750: T504 = 1'h0;
    2751: T504 = 1'h0;
    2752: T504 = 1'h0;
    2753: T504 = 1'h0;
    2754: T504 = 1'h0;
    2755: T504 = 1'h0;
    2756: T504 = 1'h0;
    2757: T504 = 1'h0;
    2758: T504 = 1'h0;
    2759: T504 = 1'h0;
    2760: T504 = 1'h0;
    2761: T504 = 1'h0;
    2762: T504 = 1'h0;
    2763: T504 = 1'h0;
    2764: T504 = 1'h0;
    2765: T504 = 1'h0;
    2766: T504 = 1'h0;
    2767: T504 = 1'h0;
    2768: T504 = 1'h0;
    2769: T504 = 1'h0;
    2770: T504 = 1'h0;
    2771: T504 = 1'h0;
    2772: T504 = 1'h0;
    2773: T504 = 1'h0;
    2774: T504 = 1'h0;
    2775: T504 = 1'h0;
    2776: T504 = 1'h0;
    2777: T504 = 1'h0;
    2778: T504 = 1'h0;
    2779: T504 = 1'h0;
    2780: T504 = 1'h0;
    2781: T504 = 1'h0;
    2782: T504 = 1'h0;
    2783: T504 = 1'h0;
    2784: T504 = 1'h0;
    2785: T504 = 1'h0;
    2786: T504 = 1'h0;
    2787: T504 = 1'h0;
    2788: T504 = 1'h0;
    2789: T504 = 1'h0;
    2790: T504 = 1'h0;
    2791: T504 = 1'h0;
    2792: T504 = 1'h0;
    2793: T504 = 1'h0;
    2794: T504 = 1'h0;
    2795: T504 = 1'h0;
    2796: T504 = 1'h0;
    2797: T504 = 1'h0;
    2798: T504 = 1'h0;
    2799: T504 = 1'h0;
    2800: T504 = 1'h0;
    2801: T504 = 1'h0;
    2802: T504 = 1'h0;
    2803: T504 = 1'h0;
    2804: T504 = 1'h0;
    2805: T504 = 1'h0;
    2806: T504 = 1'h0;
    2807: T504 = 1'h0;
    2808: T504 = 1'h0;
    2809: T504 = 1'h0;
    2810: T504 = 1'h0;
    2811: T504 = 1'h0;
    2812: T504 = 1'h0;
    2813: T504 = 1'h0;
    2814: T504 = 1'h0;
    2815: T504 = 1'h0;
    2816: T504 = 1'h0;
    2817: T504 = 1'h0;
    2818: T504 = 1'h0;
    2819: T504 = 1'h0;
    2820: T504 = 1'h0;
    2821: T504 = 1'h0;
    2822: T504 = 1'h0;
    2823: T504 = 1'h0;
    2824: T504 = 1'h0;
    2825: T504 = 1'h0;
    2826: T504 = 1'h0;
    2827: T504 = 1'h0;
    2828: T504 = 1'h0;
    2829: T504 = 1'h0;
    2830: T504 = 1'h0;
    2831: T504 = 1'h0;
    2832: T504 = 1'h0;
    2833: T504 = 1'h0;
    2834: T504 = 1'h0;
    2835: T504 = 1'h0;
    2836: T504 = 1'h0;
    2837: T504 = 1'h0;
    2838: T504 = 1'h0;
    2839: T504 = 1'h0;
    2840: T504 = 1'h0;
    2841: T504 = 1'h0;
    2842: T504 = 1'h0;
    2843: T504 = 1'h0;
    2844: T504 = 1'h0;
    2845: T504 = 1'h0;
    2846: T504 = 1'h0;
    2847: T504 = 1'h0;
    2848: T504 = 1'h0;
    2849: T504 = 1'h0;
    2850: T504 = 1'h0;
    2851: T504 = 1'h0;
    2852: T504 = 1'h0;
    2853: T504 = 1'h0;
    2854: T504 = 1'h0;
    2855: T504 = 1'h0;
    2856: T504 = 1'h0;
    2857: T504 = 1'h0;
    2858: T504 = 1'h0;
    2859: T504 = 1'h0;
    2860: T504 = 1'h0;
    2861: T504 = 1'h0;
    2862: T504 = 1'h0;
    2863: T504 = 1'h0;
    2864: T504 = 1'h0;
    2865: T504 = 1'h0;
    2866: T504 = 1'h0;
    2867: T504 = 1'h0;
    2868: T504 = 1'h0;
    2869: T504 = 1'h0;
    2870: T504 = 1'h0;
    2871: T504 = 1'h0;
    2872: T504 = 1'h0;
    2873: T504 = 1'h0;
    2874: T504 = 1'h0;
    2875: T504 = 1'h0;
    2876: T504 = 1'h0;
    2877: T504 = 1'h0;
    2878: T504 = 1'h0;
    2879: T504 = 1'h0;
    2880: T504 = 1'h0;
    2881: T504 = 1'h0;
    2882: T504 = 1'h0;
    2883: T504 = 1'h0;
    2884: T504 = 1'h0;
    2885: T504 = 1'h0;
    2886: T504 = 1'h0;
    2887: T504 = 1'h0;
    2888: T504 = 1'h0;
    2889: T504 = 1'h0;
    2890: T504 = 1'h0;
    2891: T504 = 1'h0;
    2892: T504 = 1'h0;
    2893: T504 = 1'h0;
    2894: T504 = 1'h0;
    2895: T504 = 1'h0;
    2896: T504 = 1'h0;
    2897: T504 = 1'h0;
    2898: T504 = 1'h0;
    2899: T504 = 1'h0;
    2900: T504 = 1'h0;
    2901: T504 = 1'h0;
    2902: T504 = 1'h0;
    2903: T504 = 1'h0;
    2904: T504 = 1'h0;
    2905: T504 = 1'h0;
    2906: T504 = 1'h0;
    2907: T504 = 1'h0;
    2908: T504 = 1'h0;
    2909: T504 = 1'h0;
    2910: T504 = 1'h0;
    2911: T504 = 1'h0;
    2912: T504 = 1'h0;
    2913: T504 = 1'h0;
    2914: T504 = 1'h0;
    2915: T504 = 1'h0;
    2916: T504 = 1'h0;
    2917: T504 = 1'h0;
    2918: T504 = 1'h0;
    2919: T504 = 1'h0;
    2920: T504 = 1'h0;
    2921: T504 = 1'h0;
    2922: T504 = 1'h0;
    2923: T504 = 1'h0;
    2924: T504 = 1'h0;
    2925: T504 = 1'h0;
    2926: T504 = 1'h0;
    2927: T504 = 1'h0;
    2928: T504 = 1'h0;
    2929: T504 = 1'h0;
    2930: T504 = 1'h0;
    2931: T504 = 1'h0;
    2932: T504 = 1'h0;
    2933: T504 = 1'h0;
    2934: T504 = 1'h0;
    2935: T504 = 1'h0;
    2936: T504 = 1'h0;
    2937: T504 = 1'h0;
    2938: T504 = 1'h0;
    2939: T504 = 1'h0;
    2940: T504 = 1'h0;
    2941: T504 = 1'h0;
    2942: T504 = 1'h0;
    2943: T504 = 1'h0;
    2944: T504 = 1'h0;
    2945: T504 = 1'h0;
    2946: T504 = 1'h0;
    2947: T504 = 1'h0;
    2948: T504 = 1'h0;
    2949: T504 = 1'h0;
    2950: T504 = 1'h0;
    2951: T504 = 1'h0;
    2952: T504 = 1'h0;
    2953: T504 = 1'h0;
    2954: T504 = 1'h0;
    2955: T504 = 1'h0;
    2956: T504 = 1'h0;
    2957: T504 = 1'h0;
    2958: T504 = 1'h0;
    2959: T504 = 1'h0;
    2960: T504 = 1'h0;
    2961: T504 = 1'h0;
    2962: T504 = 1'h0;
    2963: T504 = 1'h0;
    2964: T504 = 1'h0;
    2965: T504 = 1'h0;
    2966: T504 = 1'h0;
    2967: T504 = 1'h0;
    2968: T504 = 1'h0;
    2969: T504 = 1'h0;
    2970: T504 = 1'h0;
    2971: T504 = 1'h0;
    2972: T504 = 1'h0;
    2973: T504 = 1'h0;
    2974: T504 = 1'h0;
    2975: T504 = 1'h0;
    2976: T504 = 1'h0;
    2977: T504 = 1'h0;
    2978: T504 = 1'h0;
    2979: T504 = 1'h0;
    2980: T504 = 1'h0;
    2981: T504 = 1'h0;
    2982: T504 = 1'h0;
    2983: T504 = 1'h0;
    2984: T504 = 1'h0;
    2985: T504 = 1'h0;
    2986: T504 = 1'h0;
    2987: T504 = 1'h0;
    2988: T504 = 1'h0;
    2989: T504 = 1'h0;
    2990: T504 = 1'h0;
    2991: T504 = 1'h0;
    2992: T504 = 1'h0;
    2993: T504 = 1'h0;
    2994: T504 = 1'h0;
    2995: T504 = 1'h0;
    2996: T504 = 1'h0;
    2997: T504 = 1'h0;
    2998: T504 = 1'h0;
    2999: T504 = 1'h0;
    3000: T504 = 1'h0;
    3001: T504 = 1'h0;
    3002: T504 = 1'h0;
    3003: T504 = 1'h0;
    3004: T504 = 1'h0;
    3005: T504 = 1'h0;
    3006: T504 = 1'h0;
    3007: T504 = 1'h0;
    3008: T504 = 1'h0;
    3009: T504 = 1'h0;
    3010: T504 = 1'h0;
    3011: T504 = 1'h0;
    3012: T504 = 1'h0;
    3013: T504 = 1'h0;
    3014: T504 = 1'h0;
    3015: T504 = 1'h0;
    3016: T504 = 1'h0;
    3017: T504 = 1'h0;
    3018: T504 = 1'h0;
    3019: T504 = 1'h0;
    3020: T504 = 1'h0;
    3021: T504 = 1'h0;
    3022: T504 = 1'h0;
    3023: T504 = 1'h0;
    3024: T504 = 1'h0;
    3025: T504 = 1'h0;
    3026: T504 = 1'h0;
    3027: T504 = 1'h0;
    3028: T504 = 1'h0;
    3029: T504 = 1'h0;
    3030: T504 = 1'h0;
    3031: T504 = 1'h0;
    3032: T504 = 1'h0;
    3033: T504 = 1'h0;
    3034: T504 = 1'h0;
    3035: T504 = 1'h0;
    3036: T504 = 1'h0;
    3037: T504 = 1'h0;
    3038: T504 = 1'h0;
    3039: T504 = 1'h0;
    3040: T504 = 1'h0;
    3041: T504 = 1'h0;
    3042: T504 = 1'h0;
    3043: T504 = 1'h0;
    3044: T504 = 1'h0;
    3045: T504 = 1'h0;
    3046: T504 = 1'h0;
    3047: T504 = 1'h0;
    3048: T504 = 1'h0;
    3049: T504 = 1'h0;
    3050: T504 = 1'h0;
    3051: T504 = 1'h0;
    3052: T504 = 1'h0;
    3053: T504 = 1'h0;
    3054: T504 = 1'h0;
    3055: T504 = 1'h0;
    3056: T504 = 1'h0;
    3057: T504 = 1'h0;
    3058: T504 = 1'h0;
    3059: T504 = 1'h0;
    3060: T504 = 1'h0;
    3061: T504 = 1'h0;
    3062: T504 = 1'h0;
    3063: T504 = 1'h0;
    3064: T504 = 1'h0;
    3065: T504 = 1'h0;
    3066: T504 = 1'h0;
    3067: T504 = 1'h0;
    3068: T504 = 1'h0;
    3069: T504 = 1'h0;
    3070: T504 = 1'h0;
    3071: T504 = 1'h0;
    3072: T504 = 1'h1;
    3073: T504 = 1'h1;
    3074: T504 = 1'h1;
    3075: T504 = 1'h0;
    3076: T504 = 1'h0;
    3077: T504 = 1'h0;
    3078: T504 = 1'h0;
    3079: T504 = 1'h0;
    3080: T504 = 1'h0;
    3081: T504 = 1'h0;
    3082: T504 = 1'h0;
    3083: T504 = 1'h0;
    3084: T504 = 1'h0;
    3085: T504 = 1'h0;
    3086: T504 = 1'h0;
    3087: T504 = 1'h0;
    3088: T504 = 1'h0;
    3089: T504 = 1'h0;
    3090: T504 = 1'h0;
    3091: T504 = 1'h0;
    3092: T504 = 1'h0;
    3093: T504 = 1'h0;
    3094: T504 = 1'h0;
    3095: T504 = 1'h0;
    3096: T504 = 1'h0;
    3097: T504 = 1'h0;
    3098: T504 = 1'h0;
    3099: T504 = 1'h0;
    3100: T504 = 1'h0;
    3101: T504 = 1'h0;
    3102: T504 = 1'h0;
    3103: T504 = 1'h0;
    3104: T504 = 1'h0;
    3105: T504 = 1'h0;
    3106: T504 = 1'h0;
    3107: T504 = 1'h0;
    3108: T504 = 1'h0;
    3109: T504 = 1'h0;
    3110: T504 = 1'h0;
    3111: T504 = 1'h0;
    3112: T504 = 1'h0;
    3113: T504 = 1'h0;
    3114: T504 = 1'h0;
    3115: T504 = 1'h0;
    3116: T504 = 1'h0;
    3117: T504 = 1'h0;
    3118: T504 = 1'h0;
    3119: T504 = 1'h0;
    3120: T504 = 1'h0;
    3121: T504 = 1'h0;
    3122: T504 = 1'h0;
    3123: T504 = 1'h0;
    3124: T504 = 1'h0;
    3125: T504 = 1'h0;
    3126: T504 = 1'h0;
    3127: T504 = 1'h0;
    3128: T504 = 1'h0;
    3129: T504 = 1'h0;
    3130: T504 = 1'h0;
    3131: T504 = 1'h0;
    3132: T504 = 1'h0;
    3133: T504 = 1'h0;
    3134: T504 = 1'h0;
    3135: T504 = 1'h0;
    3136: T504 = 1'h0;
    3137: T504 = 1'h0;
    3138: T504 = 1'h0;
    3139: T504 = 1'h0;
    3140: T504 = 1'h0;
    3141: T504 = 1'h0;
    3142: T504 = 1'h0;
    3143: T504 = 1'h0;
    3144: T504 = 1'h0;
    3145: T504 = 1'h0;
    3146: T504 = 1'h0;
    3147: T504 = 1'h0;
    3148: T504 = 1'h0;
    3149: T504 = 1'h0;
    3150: T504 = 1'h0;
    3151: T504 = 1'h0;
    3152: T504 = 1'h0;
    3153: T504 = 1'h0;
    3154: T504 = 1'h0;
    3155: T504 = 1'h0;
    3156: T504 = 1'h0;
    3157: T504 = 1'h0;
    3158: T504 = 1'h0;
    3159: T504 = 1'h0;
    3160: T504 = 1'h0;
    3161: T504 = 1'h0;
    3162: T504 = 1'h0;
    3163: T504 = 1'h0;
    3164: T504 = 1'h0;
    3165: T504 = 1'h0;
    3166: T504 = 1'h0;
    3167: T504 = 1'h0;
    3168: T504 = 1'h0;
    3169: T504 = 1'h0;
    3170: T504 = 1'h0;
    3171: T504 = 1'h0;
    3172: T504 = 1'h0;
    3173: T504 = 1'h0;
    3174: T504 = 1'h0;
    3175: T504 = 1'h0;
    3176: T504 = 1'h0;
    3177: T504 = 1'h0;
    3178: T504 = 1'h0;
    3179: T504 = 1'h0;
    3180: T504 = 1'h0;
    3181: T504 = 1'h0;
    3182: T504 = 1'h0;
    3183: T504 = 1'h0;
    3184: T504 = 1'h0;
    3185: T504 = 1'h0;
    3186: T504 = 1'h0;
    3187: T504 = 1'h0;
    3188: T504 = 1'h0;
    3189: T504 = 1'h0;
    3190: T504 = 1'h0;
    3191: T504 = 1'h0;
    3192: T504 = 1'h0;
    3193: T504 = 1'h0;
    3194: T504 = 1'h0;
    3195: T504 = 1'h0;
    3196: T504 = 1'h0;
    3197: T504 = 1'h0;
    3198: T504 = 1'h0;
    3199: T504 = 1'h0;
    3200: T504 = 1'h0;
    3201: T504 = 1'h0;
    3202: T504 = 1'h0;
    3203: T504 = 1'h0;
    3204: T504 = 1'h0;
    3205: T504 = 1'h0;
    3206: T504 = 1'h0;
    3207: T504 = 1'h0;
    3208: T504 = 1'h0;
    3209: T504 = 1'h0;
    3210: T504 = 1'h0;
    3211: T504 = 1'h0;
    3212: T504 = 1'h0;
    3213: T504 = 1'h0;
    3214: T504 = 1'h0;
    3215: T504 = 1'h0;
    3216: T504 = 1'h0;
    3217: T504 = 1'h0;
    3218: T504 = 1'h0;
    3219: T504 = 1'h0;
    3220: T504 = 1'h0;
    3221: T504 = 1'h0;
    3222: T504 = 1'h0;
    3223: T504 = 1'h0;
    3224: T504 = 1'h0;
    3225: T504 = 1'h0;
    3226: T504 = 1'h0;
    3227: T504 = 1'h0;
    3228: T504 = 1'h0;
    3229: T504 = 1'h0;
    3230: T504 = 1'h0;
    3231: T504 = 1'h0;
    3232: T504 = 1'h0;
    3233: T504 = 1'h0;
    3234: T504 = 1'h0;
    3235: T504 = 1'h0;
    3236: T504 = 1'h0;
    3237: T504 = 1'h0;
    3238: T504 = 1'h0;
    3239: T504 = 1'h0;
    3240: T504 = 1'h0;
    3241: T504 = 1'h0;
    3242: T504 = 1'h0;
    3243: T504 = 1'h0;
    3244: T504 = 1'h0;
    3245: T504 = 1'h0;
    3246: T504 = 1'h0;
    3247: T504 = 1'h0;
    3248: T504 = 1'h0;
    3249: T504 = 1'h0;
    3250: T504 = 1'h0;
    3251: T504 = 1'h0;
    3252: T504 = 1'h0;
    3253: T504 = 1'h0;
    3254: T504 = 1'h0;
    3255: T504 = 1'h0;
    3256: T504 = 1'h0;
    3257: T504 = 1'h0;
    3258: T504 = 1'h0;
    3259: T504 = 1'h0;
    3260: T504 = 1'h0;
    3261: T504 = 1'h0;
    3262: T504 = 1'h0;
    3263: T504 = 1'h0;
    3264: T504 = 1'h1;
    3265: T504 = 1'h1;
    3266: T504 = 1'h1;
    3267: T504 = 1'h1;
    3268: T504 = 1'h1;
    3269: T504 = 1'h1;
    3270: T504 = 1'h1;
    3271: T504 = 1'h1;
    3272: T504 = 1'h1;
    3273: T504 = 1'h1;
    3274: T504 = 1'h1;
    3275: T504 = 1'h1;
    3276: T504 = 1'h1;
    3277: T504 = 1'h1;
    3278: T504 = 1'h1;
    3279: T504 = 1'h1;
    3280: T504 = 1'h0;
    3281: T504 = 1'h0;
    3282: T504 = 1'h0;
    3283: T504 = 1'h0;
    3284: T504 = 1'h0;
    3285: T504 = 1'h0;
    3286: T504 = 1'h0;
    3287: T504 = 1'h0;
    3288: T504 = 1'h0;
    3289: T504 = 1'h0;
    3290: T504 = 1'h0;
    3291: T504 = 1'h0;
    3292: T504 = 1'h0;
    3293: T504 = 1'h0;
    3294: T504 = 1'h0;
    3295: T504 = 1'h0;
    3296: T504 = 1'h0;
    3297: T504 = 1'h0;
    3298: T504 = 1'h0;
    3299: T504 = 1'h0;
    3300: T504 = 1'h0;
    3301: T504 = 1'h0;
    3302: T504 = 1'h0;
    3303: T504 = 1'h0;
    3304: T504 = 1'h0;
    3305: T504 = 1'h0;
    3306: T504 = 1'h0;
    3307: T504 = 1'h0;
    3308: T504 = 1'h0;
    3309: T504 = 1'h0;
    3310: T504 = 1'h0;
    3311: T504 = 1'h0;
    3312: T504 = 1'h0;
    3313: T504 = 1'h0;
    3314: T504 = 1'h0;
    3315: T504 = 1'h0;
    3316: T504 = 1'h0;
    3317: T504 = 1'h0;
    3318: T504 = 1'h0;
    3319: T504 = 1'h0;
    3320: T504 = 1'h0;
    3321: T504 = 1'h0;
    3322: T504 = 1'h0;
    3323: T504 = 1'h0;
    3324: T504 = 1'h0;
    3325: T504 = 1'h0;
    3326: T504 = 1'h0;
    3327: T504 = 1'h0;
    3328: T504 = 1'h0;
    3329: T504 = 1'h0;
    3330: T504 = 1'h0;
    3331: T504 = 1'h0;
    3332: T504 = 1'h0;
    3333: T504 = 1'h0;
    3334: T504 = 1'h0;
    3335: T504 = 1'h0;
    3336: T504 = 1'h0;
    3337: T504 = 1'h0;
    3338: T504 = 1'h0;
    3339: T504 = 1'h0;
    3340: T504 = 1'h0;
    3341: T504 = 1'h0;
    3342: T504 = 1'h0;
    3343: T504 = 1'h0;
    3344: T504 = 1'h0;
    3345: T504 = 1'h0;
    3346: T504 = 1'h0;
    3347: T504 = 1'h0;
    3348: T504 = 1'h0;
    3349: T504 = 1'h0;
    3350: T504 = 1'h0;
    3351: T504 = 1'h0;
    3352: T504 = 1'h0;
    3353: T504 = 1'h0;
    3354: T504 = 1'h0;
    3355: T504 = 1'h0;
    3356: T504 = 1'h0;
    3357: T504 = 1'h0;
    3358: T504 = 1'h0;
    3359: T504 = 1'h0;
    3360: T504 = 1'h0;
    3361: T504 = 1'h0;
    3362: T504 = 1'h0;
    3363: T504 = 1'h0;
    3364: T504 = 1'h0;
    3365: T504 = 1'h0;
    3366: T504 = 1'h0;
    3367: T504 = 1'h0;
    3368: T504 = 1'h0;
    3369: T504 = 1'h0;
    3370: T504 = 1'h0;
    3371: T504 = 1'h0;
    3372: T504 = 1'h0;
    3373: T504 = 1'h0;
    3374: T504 = 1'h0;
    3375: T504 = 1'h0;
    3376: T504 = 1'h0;
    3377: T504 = 1'h0;
    3378: T504 = 1'h0;
    3379: T504 = 1'h0;
    3380: T504 = 1'h0;
    3381: T504 = 1'h0;
    3382: T504 = 1'h0;
    3383: T504 = 1'h0;
    3384: T504 = 1'h0;
    3385: T504 = 1'h0;
    3386: T504 = 1'h0;
    3387: T504 = 1'h0;
    3388: T504 = 1'h0;
    3389: T504 = 1'h0;
    3390: T504 = 1'h0;
    3391: T504 = 1'h0;
    3392: T504 = 1'h0;
    3393: T504 = 1'h0;
    3394: T504 = 1'h0;
    3395: T504 = 1'h0;
    3396: T504 = 1'h0;
    3397: T504 = 1'h0;
    3398: T504 = 1'h0;
    3399: T504 = 1'h0;
    3400: T504 = 1'h0;
    3401: T504 = 1'h0;
    3402: T504 = 1'h0;
    3403: T504 = 1'h0;
    3404: T504 = 1'h0;
    3405: T504 = 1'h0;
    3406: T504 = 1'h0;
    3407: T504 = 1'h0;
    3408: T504 = 1'h0;
    3409: T504 = 1'h0;
    3410: T504 = 1'h0;
    3411: T504 = 1'h0;
    3412: T504 = 1'h0;
    3413: T504 = 1'h0;
    3414: T504 = 1'h0;
    3415: T504 = 1'h0;
    3416: T504 = 1'h0;
    3417: T504 = 1'h0;
    3418: T504 = 1'h0;
    3419: T504 = 1'h0;
    3420: T504 = 1'h0;
    3421: T504 = 1'h0;
    3422: T504 = 1'h0;
    3423: T504 = 1'h0;
    3424: T504 = 1'h0;
    3425: T504 = 1'h0;
    3426: T504 = 1'h0;
    3427: T504 = 1'h0;
    3428: T504 = 1'h0;
    3429: T504 = 1'h0;
    3430: T504 = 1'h0;
    3431: T504 = 1'h0;
    3432: T504 = 1'h0;
    3433: T504 = 1'h0;
    3434: T504 = 1'h0;
    3435: T504 = 1'h0;
    3436: T504 = 1'h0;
    3437: T504 = 1'h0;
    3438: T504 = 1'h0;
    3439: T504 = 1'h0;
    3440: T504 = 1'h0;
    3441: T504 = 1'h0;
    3442: T504 = 1'h0;
    3443: T504 = 1'h0;
    3444: T504 = 1'h0;
    3445: T504 = 1'h0;
    3446: T504 = 1'h0;
    3447: T504 = 1'h0;
    3448: T504 = 1'h0;
    3449: T504 = 1'h0;
    3450: T504 = 1'h0;
    3451: T504 = 1'h0;
    3452: T504 = 1'h0;
    3453: T504 = 1'h0;
    3454: T504 = 1'h0;
    3455: T504 = 1'h0;
    3456: T504 = 1'h0;
    3457: T504 = 1'h0;
    3458: T504 = 1'h0;
    3459: T504 = 1'h0;
    3460: T504 = 1'h0;
    3461: T504 = 1'h0;
    3462: T504 = 1'h0;
    3463: T504 = 1'h0;
    3464: T504 = 1'h0;
    3465: T504 = 1'h0;
    3466: T504 = 1'h0;
    3467: T504 = 1'h0;
    3468: T504 = 1'h0;
    3469: T504 = 1'h0;
    3470: T504 = 1'h0;
    3471: T504 = 1'h0;
    3472: T504 = 1'h0;
    3473: T504 = 1'h0;
    3474: T504 = 1'h0;
    3475: T504 = 1'h0;
    3476: T504 = 1'h0;
    3477: T504 = 1'h0;
    3478: T504 = 1'h0;
    3479: T504 = 1'h0;
    3480: T504 = 1'h0;
    3481: T504 = 1'h0;
    3482: T504 = 1'h0;
    3483: T504 = 1'h0;
    3484: T504 = 1'h0;
    3485: T504 = 1'h0;
    3486: T504 = 1'h0;
    3487: T504 = 1'h0;
    3488: T504 = 1'h0;
    3489: T504 = 1'h0;
    3490: T504 = 1'h0;
    3491: T504 = 1'h0;
    3492: T504 = 1'h0;
    3493: T504 = 1'h0;
    3494: T504 = 1'h0;
    3495: T504 = 1'h0;
    3496: T504 = 1'h0;
    3497: T504 = 1'h0;
    3498: T504 = 1'h0;
    3499: T504 = 1'h0;
    3500: T504 = 1'h0;
    3501: T504 = 1'h0;
    3502: T504 = 1'h0;
    3503: T504 = 1'h0;
    3504: T504 = 1'h0;
    3505: T504 = 1'h0;
    3506: T504 = 1'h0;
    3507: T504 = 1'h0;
    3508: T504 = 1'h0;
    3509: T504 = 1'h0;
    3510: T504 = 1'h0;
    3511: T504 = 1'h0;
    3512: T504 = 1'h0;
    3513: T504 = 1'h0;
    3514: T504 = 1'h0;
    3515: T504 = 1'h0;
    3516: T504 = 1'h0;
    3517: T504 = 1'h0;
    3518: T504 = 1'h0;
    3519: T504 = 1'h0;
    3520: T504 = 1'h0;
    3521: T504 = 1'h0;
    3522: T504 = 1'h0;
    3523: T504 = 1'h0;
    3524: T504 = 1'h0;
    3525: T504 = 1'h0;
    3526: T504 = 1'h0;
    3527: T504 = 1'h0;
    3528: T504 = 1'h0;
    3529: T504 = 1'h0;
    3530: T504 = 1'h0;
    3531: T504 = 1'h0;
    3532: T504 = 1'h0;
    3533: T504 = 1'h0;
    3534: T504 = 1'h0;
    3535: T504 = 1'h0;
    3536: T504 = 1'h0;
    3537: T504 = 1'h0;
    3538: T504 = 1'h0;
    3539: T504 = 1'h0;
    3540: T504 = 1'h0;
    3541: T504 = 1'h0;
    3542: T504 = 1'h0;
    3543: T504 = 1'h0;
    3544: T504 = 1'h0;
    3545: T504 = 1'h0;
    3546: T504 = 1'h0;
    3547: T504 = 1'h0;
    3548: T504 = 1'h0;
    3549: T504 = 1'h0;
    3550: T504 = 1'h0;
    3551: T504 = 1'h0;
    3552: T504 = 1'h0;
    3553: T504 = 1'h0;
    3554: T504 = 1'h0;
    3555: T504 = 1'h0;
    3556: T504 = 1'h0;
    3557: T504 = 1'h0;
    3558: T504 = 1'h0;
    3559: T504 = 1'h0;
    3560: T504 = 1'h0;
    3561: T504 = 1'h0;
    3562: T504 = 1'h0;
    3563: T504 = 1'h0;
    3564: T504 = 1'h0;
    3565: T504 = 1'h0;
    3566: T504 = 1'h0;
    3567: T504 = 1'h0;
    3568: T504 = 1'h0;
    3569: T504 = 1'h0;
    3570: T504 = 1'h0;
    3571: T504 = 1'h0;
    3572: T504 = 1'h0;
    3573: T504 = 1'h0;
    3574: T504 = 1'h0;
    3575: T504 = 1'h0;
    3576: T504 = 1'h0;
    3577: T504 = 1'h0;
    3578: T504 = 1'h0;
    3579: T504 = 1'h0;
    3580: T504 = 1'h0;
    3581: T504 = 1'h0;
    3582: T504 = 1'h0;
    3583: T504 = 1'h0;
    3584: T504 = 1'h0;
    3585: T504 = 1'h0;
    3586: T504 = 1'h0;
    3587: T504 = 1'h0;
    3588: T504 = 1'h0;
    3589: T504 = 1'h0;
    3590: T504 = 1'h0;
    3591: T504 = 1'h0;
    3592: T504 = 1'h0;
    3593: T504 = 1'h0;
    3594: T504 = 1'h0;
    3595: T504 = 1'h0;
    3596: T504 = 1'h0;
    3597: T504 = 1'h0;
    3598: T504 = 1'h0;
    3599: T504 = 1'h0;
    3600: T504 = 1'h0;
    3601: T504 = 1'h0;
    3602: T504 = 1'h0;
    3603: T504 = 1'h0;
    3604: T504 = 1'h0;
    3605: T504 = 1'h0;
    3606: T504 = 1'h0;
    3607: T504 = 1'h0;
    3608: T504 = 1'h0;
    3609: T504 = 1'h0;
    3610: T504 = 1'h0;
    3611: T504 = 1'h0;
    3612: T504 = 1'h0;
    3613: T504 = 1'h0;
    3614: T504 = 1'h0;
    3615: T504 = 1'h0;
    3616: T504 = 1'h0;
    3617: T504 = 1'h0;
    3618: T504 = 1'h0;
    3619: T504 = 1'h0;
    3620: T504 = 1'h0;
    3621: T504 = 1'h0;
    3622: T504 = 1'h0;
    3623: T504 = 1'h0;
    3624: T504 = 1'h0;
    3625: T504 = 1'h0;
    3626: T504 = 1'h0;
    3627: T504 = 1'h0;
    3628: T504 = 1'h0;
    3629: T504 = 1'h0;
    3630: T504 = 1'h0;
    3631: T504 = 1'h0;
    3632: T504 = 1'h0;
    3633: T504 = 1'h0;
    3634: T504 = 1'h0;
    3635: T504 = 1'h0;
    3636: T504 = 1'h0;
    3637: T504 = 1'h0;
    3638: T504 = 1'h0;
    3639: T504 = 1'h0;
    3640: T504 = 1'h0;
    3641: T504 = 1'h0;
    3642: T504 = 1'h0;
    3643: T504 = 1'h0;
    3644: T504 = 1'h0;
    3645: T504 = 1'h0;
    3646: T504 = 1'h0;
    3647: T504 = 1'h0;
    3648: T504 = 1'h0;
    3649: T504 = 1'h0;
    3650: T504 = 1'h0;
    3651: T504 = 1'h0;
    3652: T504 = 1'h0;
    3653: T504 = 1'h0;
    3654: T504 = 1'h0;
    3655: T504 = 1'h0;
    3656: T504 = 1'h0;
    3657: T504 = 1'h0;
    3658: T504 = 1'h0;
    3659: T504 = 1'h0;
    3660: T504 = 1'h0;
    3661: T504 = 1'h0;
    3662: T504 = 1'h0;
    3663: T504 = 1'h0;
    3664: T504 = 1'h0;
    3665: T504 = 1'h0;
    3666: T504 = 1'h0;
    3667: T504 = 1'h0;
    3668: T504 = 1'h0;
    3669: T504 = 1'h0;
    3670: T504 = 1'h0;
    3671: T504 = 1'h0;
    3672: T504 = 1'h0;
    3673: T504 = 1'h0;
    3674: T504 = 1'h0;
    3675: T504 = 1'h0;
    3676: T504 = 1'h0;
    3677: T504 = 1'h0;
    3678: T504 = 1'h0;
    3679: T504 = 1'h0;
    3680: T504 = 1'h0;
    3681: T504 = 1'h0;
    3682: T504 = 1'h0;
    3683: T504 = 1'h0;
    3684: T504 = 1'h0;
    3685: T504 = 1'h0;
    3686: T504 = 1'h0;
    3687: T504 = 1'h0;
    3688: T504 = 1'h0;
    3689: T504 = 1'h0;
    3690: T504 = 1'h0;
    3691: T504 = 1'h0;
    3692: T504 = 1'h0;
    3693: T504 = 1'h0;
    3694: T504 = 1'h0;
    3695: T504 = 1'h0;
    3696: T504 = 1'h0;
    3697: T504 = 1'h0;
    3698: T504 = 1'h0;
    3699: T504 = 1'h0;
    3700: T504 = 1'h0;
    3701: T504 = 1'h0;
    3702: T504 = 1'h0;
    3703: T504 = 1'h0;
    3704: T504 = 1'h0;
    3705: T504 = 1'h0;
    3706: T504 = 1'h0;
    3707: T504 = 1'h0;
    3708: T504 = 1'h0;
    3709: T504 = 1'h0;
    3710: T504 = 1'h0;
    3711: T504 = 1'h0;
    3712: T504 = 1'h0;
    3713: T504 = 1'h0;
    3714: T504 = 1'h0;
    3715: T504 = 1'h0;
    3716: T504 = 1'h0;
    3717: T504 = 1'h0;
    3718: T504 = 1'h0;
    3719: T504 = 1'h0;
    3720: T504 = 1'h0;
    3721: T504 = 1'h0;
    3722: T504 = 1'h0;
    3723: T504 = 1'h0;
    3724: T504 = 1'h0;
    3725: T504 = 1'h0;
    3726: T504 = 1'h0;
    3727: T504 = 1'h0;
    3728: T504 = 1'h0;
    3729: T504 = 1'h0;
    3730: T504 = 1'h0;
    3731: T504 = 1'h0;
    3732: T504 = 1'h0;
    3733: T504 = 1'h0;
    3734: T504 = 1'h0;
    3735: T504 = 1'h0;
    3736: T504 = 1'h0;
    3737: T504 = 1'h0;
    3738: T504 = 1'h0;
    3739: T504 = 1'h0;
    3740: T504 = 1'h0;
    3741: T504 = 1'h0;
    3742: T504 = 1'h0;
    3743: T504 = 1'h0;
    3744: T504 = 1'h0;
    3745: T504 = 1'h0;
    3746: T504 = 1'h0;
    3747: T504 = 1'h0;
    3748: T504 = 1'h0;
    3749: T504 = 1'h0;
    3750: T504 = 1'h0;
    3751: T504 = 1'h0;
    3752: T504 = 1'h0;
    3753: T504 = 1'h0;
    3754: T504 = 1'h0;
    3755: T504 = 1'h0;
    3756: T504 = 1'h0;
    3757: T504 = 1'h0;
    3758: T504 = 1'h0;
    3759: T504 = 1'h0;
    3760: T504 = 1'h0;
    3761: T504 = 1'h0;
    3762: T504 = 1'h0;
    3763: T504 = 1'h0;
    3764: T504 = 1'h0;
    3765: T504 = 1'h0;
    3766: T504 = 1'h0;
    3767: T504 = 1'h0;
    3768: T504 = 1'h0;
    3769: T504 = 1'h0;
    3770: T504 = 1'h0;
    3771: T504 = 1'h0;
    3772: T504 = 1'h0;
    3773: T504 = 1'h0;
    3774: T504 = 1'h0;
    3775: T504 = 1'h0;
    3776: T504 = 1'h0;
    3777: T504 = 1'h0;
    3778: T504 = 1'h0;
    3779: T504 = 1'h0;
    3780: T504 = 1'h0;
    3781: T504 = 1'h0;
    3782: T504 = 1'h0;
    3783: T504 = 1'h0;
    3784: T504 = 1'h0;
    3785: T504 = 1'h0;
    3786: T504 = 1'h0;
    3787: T504 = 1'h0;
    3788: T504 = 1'h0;
    3789: T504 = 1'h0;
    3790: T504 = 1'h0;
    3791: T504 = 1'h0;
    3792: T504 = 1'h0;
    3793: T504 = 1'h0;
    3794: T504 = 1'h0;
    3795: T504 = 1'h0;
    3796: T504 = 1'h0;
    3797: T504 = 1'h0;
    3798: T504 = 1'h0;
    3799: T504 = 1'h0;
    3800: T504 = 1'h0;
    3801: T504 = 1'h0;
    3802: T504 = 1'h0;
    3803: T504 = 1'h0;
    3804: T504 = 1'h0;
    3805: T504 = 1'h0;
    3806: T504 = 1'h0;
    3807: T504 = 1'h0;
    3808: T504 = 1'h0;
    3809: T504 = 1'h0;
    3810: T504 = 1'h0;
    3811: T504 = 1'h0;
    3812: T504 = 1'h0;
    3813: T504 = 1'h0;
    3814: T504 = 1'h0;
    3815: T504 = 1'h0;
    3816: T504 = 1'h0;
    3817: T504 = 1'h0;
    3818: T504 = 1'h0;
    3819: T504 = 1'h0;
    3820: T504 = 1'h0;
    3821: T504 = 1'h0;
    3822: T504 = 1'h0;
    3823: T504 = 1'h0;
    3824: T504 = 1'h0;
    3825: T504 = 1'h0;
    3826: T504 = 1'h0;
    3827: T504 = 1'h0;
    3828: T504 = 1'h0;
    3829: T504 = 1'h0;
    3830: T504 = 1'h0;
    3831: T504 = 1'h0;
    3832: T504 = 1'h0;
    3833: T504 = 1'h0;
    3834: T504 = 1'h0;
    3835: T504 = 1'h0;
    3836: T504 = 1'h0;
    3837: T504 = 1'h0;
    3838: T504 = 1'h0;
    3839: T504 = 1'h0;
    3840: T504 = 1'h0;
    3841: T504 = 1'h0;
    3842: T504 = 1'h0;
    3843: T504 = 1'h0;
    3844: T504 = 1'h0;
    3845: T504 = 1'h0;
    3846: T504 = 1'h0;
    3847: T504 = 1'h0;
    3848: T504 = 1'h0;
    3849: T504 = 1'h0;
    3850: T504 = 1'h0;
    3851: T504 = 1'h0;
    3852: T504 = 1'h0;
    3853: T504 = 1'h0;
    3854: T504 = 1'h0;
    3855: T504 = 1'h0;
    3856: T504 = 1'h0;
    3857: T504 = 1'h0;
    3858: T504 = 1'h0;
    3859: T504 = 1'h0;
    3860: T504 = 1'h0;
    3861: T504 = 1'h0;
    3862: T504 = 1'h0;
    3863: T504 = 1'h0;
    3864: T504 = 1'h0;
    3865: T504 = 1'h0;
    3866: T504 = 1'h0;
    3867: T504 = 1'h0;
    3868: T504 = 1'h0;
    3869: T504 = 1'h0;
    3870: T504 = 1'h0;
    3871: T504 = 1'h0;
    3872: T504 = 1'h0;
    3873: T504 = 1'h0;
    3874: T504 = 1'h0;
    3875: T504 = 1'h0;
    3876: T504 = 1'h0;
    3877: T504 = 1'h0;
    3878: T504 = 1'h0;
    3879: T504 = 1'h0;
    3880: T504 = 1'h0;
    3881: T504 = 1'h0;
    3882: T504 = 1'h0;
    3883: T504 = 1'h0;
    3884: T504 = 1'h0;
    3885: T504 = 1'h0;
    3886: T504 = 1'h0;
    3887: T504 = 1'h0;
    3888: T504 = 1'h0;
    3889: T504 = 1'h0;
    3890: T504 = 1'h0;
    3891: T504 = 1'h0;
    3892: T504 = 1'h0;
    3893: T504 = 1'h0;
    3894: T504 = 1'h0;
    3895: T504 = 1'h0;
    3896: T504 = 1'h0;
    3897: T504 = 1'h0;
    3898: T504 = 1'h0;
    3899: T504 = 1'h0;
    3900: T504 = 1'h0;
    3901: T504 = 1'h0;
    3902: T504 = 1'h0;
    3903: T504 = 1'h0;
    3904: T504 = 1'h0;
    3905: T504 = 1'h0;
    3906: T504 = 1'h0;
    3907: T504 = 1'h0;
    3908: T504 = 1'h0;
    3909: T504 = 1'h0;
    3910: T504 = 1'h0;
    3911: T504 = 1'h0;
    3912: T504 = 1'h0;
    3913: T504 = 1'h0;
    3914: T504 = 1'h0;
    3915: T504 = 1'h0;
    3916: T504 = 1'h0;
    3917: T504 = 1'h0;
    3918: T504 = 1'h0;
    3919: T504 = 1'h0;
    3920: T504 = 1'h0;
    3921: T504 = 1'h0;
    3922: T504 = 1'h0;
    3923: T504 = 1'h0;
    3924: T504 = 1'h0;
    3925: T504 = 1'h0;
    3926: T504 = 1'h0;
    3927: T504 = 1'h0;
    3928: T504 = 1'h0;
    3929: T504 = 1'h0;
    3930: T504 = 1'h0;
    3931: T504 = 1'h0;
    3932: T504 = 1'h0;
    3933: T504 = 1'h0;
    3934: T504 = 1'h0;
    3935: T504 = 1'h0;
    3936: T504 = 1'h0;
    3937: T504 = 1'h0;
    3938: T504 = 1'h0;
    3939: T504 = 1'h0;
    3940: T504 = 1'h0;
    3941: T504 = 1'h0;
    3942: T504 = 1'h0;
    3943: T504 = 1'h0;
    3944: T504 = 1'h0;
    3945: T504 = 1'h0;
    3946: T504 = 1'h0;
    3947: T504 = 1'h0;
    3948: T504 = 1'h0;
    3949: T504 = 1'h0;
    3950: T504 = 1'h0;
    3951: T504 = 1'h0;
    3952: T504 = 1'h0;
    3953: T504 = 1'h0;
    3954: T504 = 1'h0;
    3955: T504 = 1'h0;
    3956: T504 = 1'h0;
    3957: T504 = 1'h0;
    3958: T504 = 1'h0;
    3959: T504 = 1'h0;
    3960: T504 = 1'h0;
    3961: T504 = 1'h0;
    3962: T504 = 1'h0;
    3963: T504 = 1'h0;
    3964: T504 = 1'h0;
    3965: T504 = 1'h0;
    3966: T504 = 1'h0;
    3967: T504 = 1'h0;
    3968: T504 = 1'h0;
    3969: T504 = 1'h0;
    3970: T504 = 1'h0;
    3971: T504 = 1'h0;
    3972: T504 = 1'h0;
    3973: T504 = 1'h0;
    3974: T504 = 1'h0;
    3975: T504 = 1'h0;
    3976: T504 = 1'h0;
    3977: T504 = 1'h0;
    3978: T504 = 1'h0;
    3979: T504 = 1'h0;
    3980: T504 = 1'h0;
    3981: T504 = 1'h0;
    3982: T504 = 1'h0;
    3983: T504 = 1'h0;
    3984: T504 = 1'h0;
    3985: T504 = 1'h0;
    3986: T504 = 1'h0;
    3987: T504 = 1'h0;
    3988: T504 = 1'h0;
    3989: T504 = 1'h0;
    3990: T504 = 1'h0;
    3991: T504 = 1'h0;
    3992: T504 = 1'h0;
    3993: T504 = 1'h0;
    3994: T504 = 1'h0;
    3995: T504 = 1'h0;
    3996: T504 = 1'h0;
    3997: T504 = 1'h0;
    3998: T504 = 1'h0;
    3999: T504 = 1'h0;
    4000: T504 = 1'h0;
    4001: T504 = 1'h0;
    4002: T504 = 1'h0;
    4003: T504 = 1'h0;
    4004: T504 = 1'h0;
    4005: T504 = 1'h0;
    4006: T504 = 1'h0;
    4007: T504 = 1'h0;
    4008: T504 = 1'h0;
    4009: T504 = 1'h0;
    4010: T504 = 1'h0;
    4011: T504 = 1'h0;
    4012: T504 = 1'h0;
    4013: T504 = 1'h0;
    4014: T504 = 1'h0;
    4015: T504 = 1'h0;
    4016: T504 = 1'h0;
    4017: T504 = 1'h0;
    4018: T504 = 1'h0;
    4019: T504 = 1'h0;
    4020: T504 = 1'h0;
    4021: T504 = 1'h0;
    4022: T504 = 1'h0;
    4023: T504 = 1'h0;
    4024: T504 = 1'h0;
    4025: T504 = 1'h0;
    4026: T504 = 1'h0;
    4027: T504 = 1'h0;
    4028: T504 = 1'h0;
    4029: T504 = 1'h0;
    4030: T504 = 1'h0;
    4031: T504 = 1'h0;
    4032: T504 = 1'h0;
    4033: T504 = 1'h0;
    4034: T504 = 1'h0;
    4035: T504 = 1'h0;
    4036: T504 = 1'h0;
    4037: T504 = 1'h0;
    4038: T504 = 1'h0;
    4039: T504 = 1'h0;
    4040: T504 = 1'h0;
    4041: T504 = 1'h0;
    4042: T504 = 1'h0;
    4043: T504 = 1'h0;
    4044: T504 = 1'h0;
    4045: T504 = 1'h0;
    4046: T504 = 1'h0;
    4047: T504 = 1'h0;
    4048: T504 = 1'h0;
    4049: T504 = 1'h0;
    4050: T504 = 1'h0;
    4051: T504 = 1'h0;
    4052: T504 = 1'h0;
    4053: T504 = 1'h0;
    4054: T504 = 1'h0;
    4055: T504 = 1'h0;
    4056: T504 = 1'h0;
    4057: T504 = 1'h0;
    4058: T504 = 1'h0;
    4059: T504 = 1'h0;
    4060: T504 = 1'h0;
    4061: T504 = 1'h0;
    4062: T504 = 1'h0;
    4063: T504 = 1'h0;
    4064: T504 = 1'h0;
    4065: T504 = 1'h0;
    4066: T504 = 1'h0;
    4067: T504 = 1'h0;
    4068: T504 = 1'h0;
    4069: T504 = 1'h0;
    4070: T504 = 1'h0;
    4071: T504 = 1'h0;
    4072: T504 = 1'h0;
    4073: T504 = 1'h0;
    4074: T504 = 1'h0;
    4075: T504 = 1'h0;
    4076: T504 = 1'h0;
    4077: T504 = 1'h0;
    4078: T504 = 1'h0;
    4079: T504 = 1'h0;
    4080: T504 = 1'h0;
    4081: T504 = 1'h0;
    4082: T504 = 1'h0;
    4083: T504 = 1'h0;
    4084: T504 = 1'h0;
    4085: T504 = 1'h0;
    4086: T504 = 1'h0;
    4087: T504 = 1'h0;
    4088: T504 = 1'h0;
    4089: T504 = 1'h0;
    4090: T504 = 1'h0;
    4091: T504 = 1'h0;
    4092: T504 = 1'h0;
    4093: T504 = 1'h0;
    4094: T504 = 1'h0;
    4095: T504 = 1'h0;
    default: begin
      T504 = 1'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T504 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T506 = id_ctrl_legal ^ 1'h1;
  assign id_ctrl_legal = T507;
  assign T507 = T510 | T508;
  assign T508 = T509 == 32'h33;
  assign T509 = io_dpath_inst & 32'hfc007077;
  assign T510 = T513 | T511;
  assign T511 = T512 == 32'h4063;
  assign T512 = io_dpath_inst & 32'h407f;
  assign T513 = T516 | T514;
  assign T514 = T515 == 32'h1063;
  assign T515 = io_dpath_inst & 32'h306f;
  assign T516 = T519 | T517;
  assign T517 = T518 == 32'h23;
  assign T518 = io_dpath_inst & 32'h603f;
  assign T519 = T522 | T520;
  assign T520 = T521 == 32'he0000053;
  assign T521 = io_dpath_inst & 32'hedf0707f;
  assign T522 = T525 | T523;
  assign T523 = T524 == 32'he0000053;
  assign T524 = io_dpath_inst & 32'hfdf0607f;
  assign T525 = T528 | T526;
  assign T526 = T527 == 32'hc0000053;
  assign T527 = io_dpath_inst & 32'hedc0007f;
  assign T528 = T531 | T529;
  assign T529 = T530 == 32'h42000053;
  assign T530 = io_dpath_inst & 32'h7ff0007f;
  assign T531 = T534 | T532;
  assign T532 = T533 == 32'h40100053;
  assign T533 = io_dpath_inst & 32'h7ff0007f;
  assign T534 = T537 | T535;
  assign T535 = T536 == 32'h20000053;
  assign T536 = io_dpath_inst & 32'h7c00507f;
  assign T537 = T540 | T538;
  assign T538 = T539 == 32'h20000053;
  assign T539 = io_dpath_inst & 32'h7c00607f;
  assign T540 = T543 | T541;
  assign T541 = T542 == 32'h20000053;
  assign T542 = io_dpath_inst & 32'hf400607f;
  assign T543 = T544 | T66;
  assign T544 = T545 | T69;
  assign T545 = T548 | T546;
  assign T546 = T547 == 32'h2004033;
  assign T547 = io_dpath_inst & 32'hfe004077;
  assign T548 = T551 | T549;
  assign T549 = T550 == 32'h5033;
  assign T550 = io_dpath_inst & 32'hbe007077;
  assign T551 = T554 | T552;
  assign T552 = T553 == 32'h501b;
  assign T553 = io_dpath_inst & 32'hbe00705f;
  assign T554 = T557 | T555;
  assign T555 = T556 == 32'h5013;
  assign T556 = io_dpath_inst & 32'hbc00707f;
  assign T557 = T560 | T558;
  assign T558 = T559 == 32'h2073;
  assign T559 = io_dpath_inst & 32'h207f;
  assign T560 = T561 | T72;
  assign T561 = T564 | T562;
  assign T562 = T563 == 32'h2013;
  assign T563 = io_dpath_inst & 32'h207f;
  assign T564 = T565 | T75;
  assign T565 = T568 | T566;
  assign T566 = T567 == 32'h101b;
  assign T567 = io_dpath_inst & 32'hfe00305f;
  assign T568 = T571 | T569;
  assign T569 = T570 == 32'h1013;
  assign T570 = io_dpath_inst & 32'hfc00305f;
  assign T571 = T574 | T572;
  assign T572 = T573 == 32'h73;
  assign T573 = io_dpath_inst & 32'h7fffffff;
  assign T574 = T577 | T575;
  assign T575 = T576 == 32'h6f;
  assign T576 = io_dpath_inst & 32'h7f;
  assign T577 = T580 | T578;
  assign T578 = T579 == 32'h63;
  assign T579 = io_dpath_inst & 32'h707b;
  assign T580 = T581 | T78;
  assign T581 = T584 | T582;
  assign T582 = T583 == 32'h53;
  assign T583 = io_dpath_inst & 32'hec00007f;
  assign T584 = T587 | T585;
  assign T585 = T586 == 32'h53;
  assign T586 = io_dpath_inst & 32'hf400007f;
  assign T587 = T590 | T588;
  assign T588 = T589 == 32'h43;
  assign T589 = io_dpath_inst & 32'h4000073;
  assign T590 = T593 | T591;
  assign T591 = T592 == 32'h33;
  assign T592 = io_dpath_inst & 32'hbe007077;
  assign T593 = T596 | T594;
  assign T594 = T595 == 32'h33;
  assign T595 = io_dpath_inst & 32'hfc00007f;
  assign T596 = T599 | T597;
  assign T597 = T598 == 32'h17;
  assign T598 = io_dpath_inst & 32'h5f;
  assign T599 = T602 | T600;
  assign T600 = T601 == 32'h13;
  assign T601 = io_dpath_inst & 32'h7077;
  assign T602 = T605 | T603;
  assign T603 = T604 == 32'hf;
  assign T604 = io_dpath_inst & 32'h607f;
  assign T605 = T84 | T606;
  assign T606 = T607 == 32'h3;
  assign T607 = io_dpath_inst & 32'h106f;
  assign T608 = T609 | io_imem_resp_bits_xcpt_if;
  assign T609 = ctrl_draind | io_imem_resp_bits_xcpt_ma;
  assign T611 = T612 & io_imem_resp_valid;
  assign T612 = ctrl_draind & T613;
  assign T613 = take_pc ^ 1'h1;
  assign T615 = dcache_kill_mem | take_pc_wb;
  assign dcache_kill_mem = T616 & io_dmem_replay_next_valid;
  assign T616 = mem_reg_valid & mem_ctrl_wxd;
  assign T617 = ctrl_killm ^ 1'h1;
  assign replay_wb_common = T618 | io_dpath_csr_replay;
  assign T618 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T619 = replay_mem & T620;
  assign T620 = take_pc_wb ^ 1'h1;
  assign replay_mem = T621 | fpu_kill_mem;
  assign T621 = dcache_kill_mem | mem_reg_replay;
  assign T622 = T623 & replay_ex;
  assign T623 = take_pc ^ 1'h1;
  assign mem_xcpt = T626 | T624;
  assign T624 = T625 & io_dmem_xcpt_pf_ld;
  assign T625 = mem_reg_valid & mem_ctrl_mem;
  assign T626 = T629 | T627;
  assign T627 = T628 & io_dmem_xcpt_pf_st;
  assign T628 = mem_reg_valid & mem_ctrl_mem;
  assign T629 = T632 | T630;
  assign T630 = T631 & io_dmem_xcpt_ma_ld;
  assign T631 = mem_reg_valid & mem_ctrl_mem;
  assign T632 = T635 | T633;
  assign T633 = T634 & io_dmem_xcpt_ma_st;
  assign T634 = mem_reg_valid & mem_ctrl_mem;
  assign T635 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T636 = T637 & ex_reg_xcpt_interrupt;
  assign T637 = take_pc ^ 1'h1;
//  assign io_rocc_pptw_sret = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_s = {1{$random}};
//  assign io_rocc_pptw_status_ps = {1{$random}};
//  assign io_rocc_pptw_status_ei = {1{$random}};
//  assign io_rocc_pptw_status_pei = {1{$random}};
//  assign io_rocc_pptw_status_ef = {1{$random}};
//  assign io_rocc_pptw_status_u64 = {1{$random}};
//  assign io_rocc_pptw_status_s64 = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_er = {1{$random}};
//  assign io_rocc_pptw_status_zero = {1{$random}};
//  assign io_rocc_pptw_status_im = {1{$random}};
//  assign io_rocc_pptw_status_ip = {1{$random}};
//  assign io_rocc_pptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_pptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_sret = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_s = {1{$random}};
//  assign io_rocc_dptw_status_ps = {1{$random}};
//  assign io_rocc_dptw_status_ei = {1{$random}};
//  assign io_rocc_dptw_status_pei = {1{$random}};
//  assign io_rocc_dptw_status_ef = {1{$random}};
//  assign io_rocc_dptw_status_u64 = {1{$random}};
//  assign io_rocc_dptw_status_s64 = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_er = {1{$random}};
//  assign io_rocc_dptw_status_zero = {1{$random}};
//  assign io_rocc_dptw_status_im = {1{$random}};
//  assign io_rocc_dptw_status_ip = {1{$random}};
//  assign io_rocc_dptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_dptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_sret = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_s = {1{$random}};
//  assign io_rocc_iptw_status_ps = {1{$random}};
//  assign io_rocc_iptw_status_ei = {1{$random}};
//  assign io_rocc_iptw_status_pei = {1{$random}};
//  assign io_rocc_iptw_status_ef = {1{$random}};
//  assign io_rocc_iptw_status_u64 = {1{$random}};
//  assign io_rocc_iptw_status_s64 = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_er = {1{$random}};
//  assign io_rocc_iptw_status_zero = {1{$random}};
//  assign io_rocc_iptw_status_im = {1{$random}};
//  assign io_rocc_iptw_status_ip = {1{$random}};
//  assign io_rocc_iptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_iptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_release_ready = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_p_type = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_addr = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_probe_valid = {1{$random}};
//  assign io_rocc_dmem_finish_ready = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_dmem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_grant_valid = {1{$random}};
//  assign io_rocc_dmem_acquire_ready = {1{$random}};
//  assign io_rocc_imem_finish_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_imem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_imem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
  assign io_rocc_s = io_dpath_status_s;
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_ptw_req_bits = {1{$random}};
//  assign io_rocc_mem_ptw_req_valid = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_data_subword = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_rocc_cmd_bits_rs2 = {2{$random}};
//  assign io_rocc_cmd_bits_rs1 = {2{$random}};
//  assign io_rocc_cmd_bits_inst_opcode = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_funct = {1{$random}};
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = T639 & T638;
  assign T638 = replay_wb_common ^ 1'h1;
  assign T639 = wb_reg_valid & wb_ctrl_rocc;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T640;
  assign T640 = T641 & id_ctrl_fp;
  assign T641 = ctrl_killd ^ 1'h1;
//  assign io_dmem_ptw_sret = {1{$random}};
//  assign io_dmem_ptw_invalidate = {1{$random}};
//  assign io_dmem_ptw_status_s = {1{$random}};
//  assign io_dmem_ptw_status_ps = {1{$random}};
//  assign io_dmem_ptw_status_ei = {1{$random}};
//  assign io_dmem_ptw_status_pei = {1{$random}};
//  assign io_dmem_ptw_status_ef = {1{$random}};
//  assign io_dmem_ptw_status_u64 = {1{$random}};
//  assign io_dmem_ptw_status_s64 = {1{$random}};
//  assign io_dmem_ptw_status_vm = {1{$random}};
//  assign io_dmem_ptw_status_er = {1{$random}};
//  assign io_dmem_ptw_status_zero = {1{$random}};
//  assign io_dmem_ptw_status_im = {1{$random}};
//  assign io_dmem_ptw_status_ip = {1{$random}};
//  assign io_dmem_ptw_resp_bits_perm = {1{$random}};
//  assign io_dmem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_dmem_ptw_resp_bits_error = {1{$random}};
//  assign io_dmem_ptw_resp_valid = {1{$random}};
//  assign io_dmem_ptw_req_ready = {1{$random}};
//  assign io_dmem_req_bits_data = {2{$random}};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
//  assign io_dmem_req_bits_tag = {1{$random}};
//  assign io_dmem_req_bits_addr = {2{$random}};
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_kill = T642;
  assign T642 = killm_common | mem_xcpt;
  assign io_dmem_req_valid = T643;
  assign T643 = ex_reg_valid & ex_ctrl_mem;
  assign io_imem_invalidate = T644;
  assign T644 = wb_reg_valid & wb_ctrl_fence_i;
  assign T645 = T452 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign T646 = T451 ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign T647 = T11 ? id_ctrl_fence_i : ex_ctrl_fence_i;
//  assign io_imem_ptw_sret = {1{$random}};
//  assign io_imem_ptw_invalidate = {1{$random}};
//  assign io_imem_ptw_status_s = {1{$random}};
//  assign io_imem_ptw_status_ps = {1{$random}};
//  assign io_imem_ptw_status_ei = {1{$random}};
//  assign io_imem_ptw_status_pei = {1{$random}};
//  assign io_imem_ptw_status_ef = {1{$random}};
//  assign io_imem_ptw_status_u64 = {1{$random}};
//  assign io_imem_ptw_status_s64 = {1{$random}};
//  assign io_imem_ptw_status_vm = {1{$random}};
//  assign io_imem_ptw_status_er = {1{$random}};
//  assign io_imem_ptw_status_zero = {1{$random}};
//  assign io_imem_ptw_status_im = {1{$random}};
//  assign io_imem_ptw_status_ip = {1{$random}};
//  assign io_imem_ptw_resp_bits_perm = {1{$random}};
//  assign io_imem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_imem_ptw_resp_bits_error = {1{$random}};
//  assign io_imem_ptw_resp_valid = {1{$random}};
//  assign io_imem_ptw_req_ready = {1{$random}};
  assign io_imem_ras_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T648 = T651 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T649 = T650 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T650 = T11 & io_imem_btb_resp_valid;
  assign T651 = T451 & ex_reg_btb_hit;
  assign T652 = T11 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T653 = T651 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T654 = T650 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T655 = T651 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T656 = T650 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_ras_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T657 = T651 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T658 = T650 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_ras_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign T659 = T651 ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign T660 = T650 ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign io_imem_ras_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign T661 = T651 ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign T662 = T650 ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign io_imem_ras_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T663 = T651 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T664 = T650 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_ras_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T665 = T451 ? ex_reg_btb_hit : mem_reg_btb_hit;
//  assign io_imem_ras_update_bits_returnAddr = {2{$random}};
  assign io_imem_ras_update_bits_isReturn = T666;
  assign T666 = mem_ctrl_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_ras_update_bits_isCall = T667;
  assign T667 = mem_ctrl_wxd & T668;
  assign T668 = io_dpath_mem_waddr[1'h0:1'h0];
  assign io_imem_ras_update_valid = T669;
  assign T669 = io_imem_btb_update_bits_isJump & T670;
  assign T670 = take_pc_wb ^ 1'h1;
  assign io_imem_bht_update_bits_mispredict = io_dpath_mem_misprediction;
  assign io_imem_bht_update_bits_taken = io_dpath_mem_br_taken;
//  assign io_imem_bht_update_bits_pc = {2{$random}};
  assign io_imem_bht_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_bht_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_bht_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_bht_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_bht_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_bht_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_bht_update_valid = T671;
  assign T671 = T673 & T672;
  assign T672 = take_pc_wb ^ 1'h1;
  assign T673 = mem_reg_valid & mem_ctrl_branch;
//  assign io_imem_btb_update_bits_br_pc = {2{$random}};
  assign io_imem_btb_update_bits_isReturn = T674;
  assign T674 = mem_ctrl_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_btb_update_bits_isJump = T675;
  assign T675 = mem_ctrl_jal | mem_ctrl_jalr;
//  assign io_imem_btb_update_bits_taken = {1{$random}};
//  assign io_imem_btb_update_bits_target = {2{$random}};
//  assign io_imem_btb_update_bits_pc = {2{$random}};
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T676;
  assign T676 = T678 & T677;
  assign T677 = take_pc_wb ^ 1'h1;
  assign T678 = T682 & T679;
  assign T679 = T680 | mem_ctrl_jal;
  assign T680 = T681 | mem_ctrl_jalr;
  assign T681 = mem_ctrl_branch & io_dpath_mem_br_taken;
  assign T682 = mem_reg_valid & io_dpath_mem_misprediction;
  assign io_imem_resp_ready = T683;
  assign T683 = T684 | ctrl_draind;
  assign T684 = ctrl_stalld ^ 1'h1;
//  assign io_imem_req_bits_pc = {2{$random}};
  assign io_imem_req_valid = take_pc;
  assign io_dpath_badvaddr_wen = wb_reg_xcpt;
  assign io_dpath_cause = wb_reg_cause;
  assign T685 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T635 ? mem_reg_cause : T908;
  assign T908 = {60'h0, T686};
  assign T686 = T633 ? 4'h9 : T687;
  assign T687 = T630 ? 4'h8 : T688;
  assign T688 = T627 ? 4'hb : 4'ha;
  assign T689 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T461 ? ex_reg_cause : 64'h2;
  assign T690 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = ctrl_draind ? id_interrupt_cause : T909;
  assign T909 = {60'h0, T691};
  assign T691 = io_imem_resp_bits_xcpt_ma ? 4'h0 : T692;
  assign T692 = io_imem_resp_bits_xcpt_if ? 4'h1 : T693;
  assign T693 = T502 ? 4'h2 : T694;
  assign T694 = id_csr_privileged ? 4'h3 : T695;
  assign T695 = T476 ? 4'h3 : T696;
  assign T696 = T470 ? 4'h4 : T697;
  assign T697 = id_ctrl_scall ? 4'h6 : 4'hc;
  assign id_interrupt_cause = T40 ? 64'h8000000000000000 : T698;
  assign T698 = T37 ? 64'h8000000000000001 : T699;
  assign T699 = T33 ? 64'h8000000000000002 : T700;
  assign T700 = T29 ? 64'h8000000000000003 : T701;
  assign T701 = T25 ? 64'h8000000000000004 : T702;
  assign T702 = T21 ? 64'h8000000000000005 : T703;
  assign T703 = T17 ? 64'h8000000000000006 : 64'h8000000000000007;
  assign io_dpath_exception = wb_reg_xcpt;
  assign io_dpath_retire = T704;
  assign T704 = wb_reg_valid & T705;
  assign T705 = replay_wb ^ 1'h1;
  assign io_dpath_ll_ready = T706;
  assign T706 = T707 ^ 1'h1;
  assign T707 = wb_reg_valid & wb_ctrl_wxd;
  assign io_dpath_bypass_src_0 = T708;
  assign T708 = T719 ? 2'h0 : T709;
  assign T709 = T716 ? 2'h1 : T710;
  assign T710 = T711 ? 2'h2 : 2'h3;
  assign T711 = T713 & T712;
  assign T712 = io_dpath_mem_waddr == id_raddr1;
  assign T713 = T715 & T714;
  assign T714 = mem_ctrl_mem ^ 1'h1;
  assign T715 = mem_reg_valid & mem_ctrl_wxd;
  assign T716 = T718 & T717;
  assign T717 = io_dpath_ex_waddr == id_raddr1;
  assign T718 = ex_reg_valid & ex_ctrl_wxd;
  assign T719 = 5'h0 == id_raddr1;
  assign io_dpath_bypass_src_1 = T720;
  assign T720 = T727 ? 2'h0 : T721;
  assign T721 = T725 ? 2'h1 : T722;
  assign T722 = T723 ? 2'h2 : 2'h3;
  assign T723 = T713 & T724;
  assign T724 = io_dpath_mem_waddr == id_raddr2;
  assign T725 = T718 & T726;
  assign T726 = io_dpath_ex_waddr == id_raddr2;
  assign T727 = 5'h0 == id_raddr2;
  assign io_dpath_bypass_0 = T728;
  assign T728 = T732 | T729;
  assign T729 = T731 & T730;
  assign T730 = io_dpath_mem_waddr == id_raddr1;
  assign T731 = mem_reg_valid & mem_ctrl_wxd;
  assign T732 = T733 | T711;
  assign T733 = T719 | T716;
  assign io_dpath_bypass_1 = T734;
  assign T734 = T737 | T735;
  assign T735 = T731 & T736;
  assign T736 = io_dpath_mem_waddr == id_raddr2;
  assign T737 = T738 | T723;
  assign T738 = T727 | T725;
  assign io_dpath_wb_wen = T739;
  assign T739 = io_dpath_retire & wb_ctrl_wxd;
  assign io_dpath_ex_valid = ex_reg_valid;
  assign io_dpath_sret = T740;
  assign T740 = T742 & T741;
  assign T741 = replay_wb ^ 1'h1;
  assign T742 = wb_reg_valid & wb_ctrl_sret;
  assign T743 = T452 ? mem_ctrl_sret : wb_ctrl_sret;
  assign T744 = T451 ? ex_ctrl_sret : mem_ctrl_sret;
  assign T745 = T11 ? id_ctrl_sret : ex_ctrl_sret;
  assign io_dpath_csr = T910;
  assign T910 = {1'h0, T746};
  assign T746 = wb_reg_valid ? wb_ctrl_csr : 2'h0;
  assign T747 = T452 ? mem_ctrl_csr : wb_ctrl_csr;
  assign io_dpath_mem_ctrl_amo = mem_ctrl_amo;
  assign T748 = T451 ? ex_ctrl_amo : mem_ctrl_amo;
  assign T749 = T11 ? id_ctrl_amo : ex_ctrl_amo;
  assign io_dpath_mem_ctrl_fence = mem_ctrl_fence;
  assign T750 = T451 ? ex_ctrl_fence : mem_ctrl_fence;
  assign T751 = T11 ? id_ctrl_fence : ex_ctrl_fence;
  assign io_dpath_mem_ctrl_scall = mem_ctrl_scall;
  assign T752 = T451 ? ex_ctrl_scall : mem_ctrl_scall;
  assign T753 = T11 ? id_ctrl_scall : ex_ctrl_scall;
  assign io_dpath_mem_ctrl_sret = mem_ctrl_sret;
  assign io_dpath_mem_ctrl_fence_i = mem_ctrl_fence_i;
  assign io_dpath_mem_ctrl_csr = mem_ctrl_csr;
  assign io_dpath_mem_ctrl_wxd = mem_ctrl_wxd;
  assign io_dpath_mem_ctrl_div = mem_ctrl_div;
  assign io_dpath_mem_ctrl_wfd = mem_ctrl_wfd;
  assign io_dpath_mem_ctrl_rfs3 = mem_ctrl_rfs3;
  assign T754 = T451 ? ex_ctrl_rfs3 : mem_ctrl_rfs3;
  assign T755 = T11 ? id_ctrl_rfs3 : ex_ctrl_rfs3;
  assign id_ctrl_rfs3 = T129;
  assign io_dpath_mem_ctrl_rfs2 = mem_ctrl_rfs2;
  assign T756 = T451 ? ex_ctrl_rfs2 : mem_ctrl_rfs2;
  assign T757 = T11 ? id_ctrl_rfs2 : ex_ctrl_rfs2;
  assign id_ctrl_rfs2 = T758;
  assign T758 = T759 | T129;
  assign T759 = T762 | T760;
  assign T760 = T761 == 32'h40;
  assign T761 = io_dpath_inst & 32'h40000064;
  assign T762 = T763 == 32'h24;
  assign T763 = io_dpath_inst & 32'h7c;
  assign io_dpath_mem_ctrl_rfs1 = mem_ctrl_rfs1;
  assign T764 = T451 ? ex_ctrl_rfs1 : mem_ctrl_rfs1;
  assign T765 = T11 ? id_ctrl_rfs1 : ex_ctrl_rfs1;
  assign id_ctrl_rfs1 = T766;
  assign T766 = T767 | T132;
  assign T767 = T768 | T129;
  assign T768 = T769 == 32'h40;
  assign T769 = io_dpath_inst & 32'h10000064;
  assign io_dpath_mem_ctrl_mem_type = mem_ctrl_mem_type;
  assign T770 = T451 ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign io_dpath_mem_ctrl_mem_cmd = mem_ctrl_mem_cmd;
  assign T771 = T451 ? ex_ctrl_mem_cmd : mem_ctrl_mem_cmd;
  assign io_dpath_mem_ctrl_mem = mem_ctrl_mem;
  assign io_dpath_mem_ctrl_alu_fn = mem_ctrl_alu_fn;
  assign T772 = T451 ? ex_ctrl_alu_fn : mem_ctrl_alu_fn;
  assign T773 = T11 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign id_ctrl_alu_fn = T774;
  assign T774 = {T810, T775};
  assign T775 = {T799, T776};
  assign T776 = {T785, T777};
  assign T777 = T780 | T778;
  assign T778 = T779 == 32'h7000;
  assign T779 = io_dpath_inst & 32'h7044;
  assign T780 = T783 | T781;
  assign T781 = T782 == 32'h1040;
  assign T782 = io_dpath_inst & 32'h1058;
  assign T783 = T784 == 32'h1010;
  assign T784 = io_dpath_inst & 32'h3054;
  assign T785 = T788 | T786;
  assign T786 = T787 == 32'h40001010;
  assign T787 = io_dpath_inst & 32'h40001054;
  assign T788 = T791 | T789;
  assign T789 = T790 == 32'h40000030;
  assign T790 = io_dpath_inst & 32'h40003034;
  assign T791 = T794 | T792;
  assign T792 = T793 == 32'h6010;
  assign T793 = io_dpath_inst & 32'h6054;
  assign T794 = T797 | T795;
  assign T795 = T796 == 32'h3010;
  assign T796 = io_dpath_inst & 32'h3054;
  assign T797 = T798 == 32'h2040;
  assign T798 = io_dpath_inst & 32'h2058;
  assign T799 = T802 | T800;
  assign T800 = T801 == 32'h4040;
  assign T801 = io_dpath_inst & 32'h4058;
  assign T802 = T805 | T803;
  assign T803 = T804 == 32'h4010;
  assign T804 = io_dpath_inst & 32'h5054;
  assign T805 = T808 | T806;
  assign T806 = T807 == 32'h4010;
  assign T807 = io_dpath_inst & 32'h40004054;
  assign T808 = T809 == 32'h2010;
  assign T809 = io_dpath_inst & 32'h2054;
  assign T810 = T813 | T811;
  assign T811 = T812 == 32'h40001010;
  assign T812 = io_dpath_inst & 32'h40003054;
  assign T813 = T814 | T789;
  assign T814 = T817 | T815;
  assign T815 = T816 == 32'h2010;
  assign T816 = io_dpath_inst & 32'h6054;
  assign T817 = T818 == 32'h40;
  assign T818 = io_dpath_inst & 32'h54;
  assign io_dpath_mem_ctrl_alu_dw = mem_ctrl_alu_dw;
  assign T819 = T451 ? ex_ctrl_alu_dw : mem_ctrl_alu_dw;
  assign T820 = T11 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign id_ctrl_alu_dw = T821;
  assign T821 = T824 | T822;
  assign T822 = T823 == 32'h0;
  assign T823 = io_dpath_inst & 32'h8;
  assign T824 = T825 == 32'h0;
  assign T825 = io_dpath_inst & 32'h10;
  assign io_dpath_mem_ctrl_sel_imm = mem_ctrl_sel_imm;
  assign T826 = T451 ? ex_ctrl_sel_imm : mem_ctrl_sel_imm;
  assign T827 = T11 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign id_ctrl_sel_imm = T828;
  assign T828 = {T838, T829};
  assign T829 = {T835, T830};
  assign T830 = T833 | T831;
  assign T831 = T832 == 32'h40;
  assign T832 = io_dpath_inst & 32'h44;
  assign T833 = T834 == 32'h8;
  assign T834 = io_dpath_inst & 32'h18;
  assign T835 = T833 | T836;
  assign T836 = T837 == 32'h14;
  assign T837 = io_dpath_inst & 32'h54;
  assign T838 = T841 | T839;
  assign T839 = T840 == 32'h40;
  assign T840 = io_dpath_inst & 32'h1060;
  assign T841 = T844 | T842;
  assign T842 = T843 == 32'h10;
  assign T843 = io_dpath_inst & 32'h14;
  assign T844 = T847 | T845;
  assign T845 = T846 == 32'h4;
  assign T846 = io_dpath_inst & 32'h201c;
  assign T847 = T848 == 32'h0;
  assign T848 = io_dpath_inst & 32'h30;
  assign io_dpath_mem_ctrl_sel_alu1 = mem_ctrl_sel_alu1;
  assign T849 = T451 ? ex_ctrl_sel_alu1 : mem_ctrl_sel_alu1;
  assign T850 = T11 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign id_ctrl_sel_alu1 = T851;
  assign T851 = {T864, T852};
  assign T852 = T855 | T853;
  assign T853 = T854 == 32'h40;
  assign T854 = io_dpath_inst & 32'h60;
  assign T855 = T858 | T856;
  assign T856 = T857 == 32'h0;
  assign T857 = io_dpath_inst & 32'h18;
  assign T858 = T859 | T278;
  assign T859 = T862 | T860;
  assign T860 = T861 == 32'h0;
  assign T861 = io_dpath_inst & 32'h50;
  assign T862 = T863 == 32'h0;
  assign T863 = io_dpath_inst & 32'h4004;
  assign T864 = T867 | T865;
  assign T865 = T866 == 32'h48;
  assign T866 = io_dpath_inst & 32'h48;
  assign T867 = T868 == 32'h14;
  assign T868 = io_dpath_inst & 32'h74;
  assign io_dpath_mem_ctrl_sel_alu2 = mem_ctrl_sel_alu2;
  assign T869 = T451 ? ex_ctrl_sel_alu2 : mem_ctrl_sel_alu2;
  assign T870 = T11 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign id_ctrl_sel_alu2 = T871;
  assign T871 = {T884, T872};
  assign T872 = T875 | T873;
  assign T873 = T874 == 32'h4050;
  assign T874 = io_dpath_inst & 32'h4050;
  assign T875 = T876 | T865;
  assign T876 = T879 | T877;
  assign T877 = T878 == 32'h4;
  assign T878 = io_dpath_inst & 32'hc;
  assign T879 = T882 | T880;
  assign T880 = T881 == 32'h0;
  assign T881 = io_dpath_inst & 32'h20;
  assign T882 = T883 == 32'h0;
  assign T883 = io_dpath_inst & 32'h58;
  assign T884 = T887 | T885;
  assign T885 = T886 == 32'h4000;
  assign T886 = io_dpath_inst & 32'h4008;
  assign T887 = T888 | T856;
  assign T888 = T889 | T880;
  assign T889 = T890 | T278;
  assign T890 = T891 == 32'h0;
  assign T891 = io_dpath_inst & 32'h48;
  assign io_dpath_mem_ctrl_rxs1 = mem_ctrl_rxs1;
  assign T892 = T451 ? ex_ctrl_rxs1 : mem_ctrl_rxs1;
  assign T893 = T11 ? id_ctrl_rxs1 : ex_ctrl_rxs1;
  assign io_dpath_mem_ctrl_rxs2 = mem_ctrl_rxs2;
  assign T894 = T451 ? ex_ctrl_rxs2 : mem_ctrl_rxs2;
  assign T895 = T11 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign io_dpath_mem_ctrl_jalr = mem_ctrl_jalr;
  assign io_dpath_mem_ctrl_jal = mem_ctrl_jal;
  assign io_dpath_mem_ctrl_branch = mem_ctrl_branch;
  assign io_dpath_mem_ctrl_rocc = mem_ctrl_rocc;
  assign io_dpath_mem_ctrl_fp = mem_ctrl_fp;
  assign io_dpath_mem_ctrl_legal = mem_ctrl_legal;
  assign T896 = T451 ? ex_ctrl_legal : mem_ctrl_legal;
  assign T897 = T11 ? id_ctrl_legal : ex_ctrl_legal;
  assign io_dpath_ex_ctrl_amo = ex_ctrl_amo;
  assign io_dpath_ex_ctrl_fence = ex_ctrl_fence;
  assign io_dpath_ex_ctrl_scall = ex_ctrl_scall;
  assign io_dpath_ex_ctrl_sret = ex_ctrl_sret;
  assign io_dpath_ex_ctrl_fence_i = ex_ctrl_fence_i;
  assign io_dpath_ex_ctrl_csr = ex_ctrl_csr;
  assign io_dpath_ex_ctrl_wxd = ex_ctrl_wxd;
  assign io_dpath_ex_ctrl_div = ex_ctrl_div;
  assign io_dpath_ex_ctrl_wfd = ex_ctrl_wfd;
  assign io_dpath_ex_ctrl_rfs3 = ex_ctrl_rfs3;
  assign io_dpath_ex_ctrl_rfs2 = ex_ctrl_rfs2;
  assign io_dpath_ex_ctrl_rfs1 = ex_ctrl_rfs1;
  assign io_dpath_ex_ctrl_mem_type = ex_ctrl_mem_type;
  assign io_dpath_ex_ctrl_mem_cmd = ex_ctrl_mem_cmd;
  assign io_dpath_ex_ctrl_mem = ex_ctrl_mem;
  assign io_dpath_ex_ctrl_alu_fn = ex_ctrl_alu_fn;
  assign io_dpath_ex_ctrl_alu_dw = ex_ctrl_alu_dw;
  assign io_dpath_ex_ctrl_sel_imm = ex_ctrl_sel_imm;
  assign io_dpath_ex_ctrl_sel_alu1 = ex_ctrl_sel_alu1;
  assign io_dpath_ex_ctrl_sel_alu2 = ex_ctrl_sel_alu2;
  assign io_dpath_ex_ctrl_rxs1 = ex_ctrl_rxs1;
  assign io_dpath_ex_ctrl_rxs2 = ex_ctrl_rxs2;
  assign io_dpath_ex_ctrl_jalr = ex_ctrl_jalr;
  assign io_dpath_ex_ctrl_jal = ex_ctrl_jal;
  assign io_dpath_ex_ctrl_branch = ex_ctrl_branch;
  assign io_dpath_ex_ctrl_rocc = ex_ctrl_rocc;
  assign io_dpath_ex_ctrl_fp = ex_ctrl_fp;
  assign io_dpath_ex_ctrl_legal = ex_ctrl_legal;
  assign io_dpath_ren_0 = id_ctrl_rxs1;
  assign io_dpath_ren_1 = id_ctrl_rxs2;
  assign io_dpath_killm = killm_common;
  assign io_dpath_killd = T898;
  assign T898 = take_pc | T899;
  assign T899 = ctrl_stalld & T900;
  assign T900 = ctrl_draind ^ 1'h1;
  assign io_dpath_sel_pc = T911;
  assign T911 = {1'h0, T901};
  assign T901 = wb_reg_xcpt ? 2'h3 : T902;
  assign T902 = replay_wb ? 2'h2 : T903;
  assign T903 = T904 ? 2'h3 : 2'h1;
  assign T904 = wb_reg_valid & wb_ctrl_sret;

  always @(posedge clk) begin
    wb_reg_xcpt <= T1;
    if(T452) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if(T451) begin
      mem_ctrl_rocc <= ex_ctrl_rocc;
    end
    if(T11) begin
      ex_ctrl_rocc <= id_ctrl_rocc;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T88;
    end
    if(reset) begin
      R112 <= 32'h0;
    end else if(T149) begin
      R112 <= T145;
    end else if(T144) begin
      R112 <= T140;
    end else if(T119) begin
      R112 <= T116;
    end
    if(T452) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if(T451) begin
      mem_ctrl_wfd <= ex_ctrl_wfd;
    end
    if(T11) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if(T452) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if(T451) begin
      mem_ctrl_mem <= ex_ctrl_mem;
    end
    if(T11) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    if(reset) begin
      R194 <= 32'h0;
    end else if(T207) begin
      R194 <= T197;
    end else if(io_dpath_ll_wen) begin
      R194 <= T190;
    end
    if(T452) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if(T451) begin
      mem_ctrl_div <= ex_ctrl_div;
    end
    if(T11) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if(T452) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if(T451) begin
      mem_ctrl_wxd <= ex_ctrl_wxd;
    end
    if(T11) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if(T451) begin
      mem_ctrl_fp <= ex_ctrl_fp;
    end
    if(T11) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    if(T451) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T11) begin
      ex_ctrl_mem_type <= id_ctrl_mem_type;
    end
    if(T11) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if(T451) begin
      mem_ctrl_csr <= ex_ctrl_csr;
    end
    if(T11) begin
      ex_ctrl_csr <= id_ctrl_csr;
    end
    mem_reg_valid <= T391;
    ex_reg_valid <= T394;
    if(T11) begin
      ex_reg_load_use <= id_load_use;
    end
    if(T451) begin
      mem_reg_flush_pipe <= ex_reg_flush_pipe;
    end
    if(T11) begin
      ex_reg_flush_pipe <= T407;
    end
    if(T451) begin
      mem_ctrl_jal <= ex_ctrl_jal;
    end
    if(T11) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if(T451) begin
      mem_ctrl_jalr <= ex_ctrl_jalr;
    end
    if(T11) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if(T451) begin
      mem_ctrl_branch <= ex_ctrl_branch;
    end
    if(T11) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if(T451) begin
      mem_reg_xcpt <= ex_xcpt;
    end else begin
      mem_reg_xcpt <= T459;
    end
    if(T11) begin
      ex_reg_xcpt <= id_xcpt;
    end else begin
      ex_reg_xcpt <= T463;
    end
    ex_reg_xcpt_interrupt <= T611;
    wb_reg_valid <= T617;
    wb_reg_replay <= T619;
    mem_reg_replay <= T622;
    mem_reg_xcpt_interrupt <= T636;
    if(T452) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if(T451) begin
      mem_ctrl_fence_i <= ex_ctrl_fence_i;
    end
    if(T11) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if(T651) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T650) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(T11) begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T651) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T650) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T651) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T650) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T651) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T650) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T651) begin
      mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
    end
    if(T650) begin
      ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
    end
    if(T651) begin
      mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
    end
    if(T650) begin
      ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
    end
    if(T651) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T650) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T451) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(T452) begin
      wb_ctrl_sret <= mem_ctrl_sret;
    end
    if(T451) begin
      mem_ctrl_sret <= ex_ctrl_sret;
    end
    if(T11) begin
      ex_ctrl_sret <= id_ctrl_sret;
    end
    if(T452) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if(T451) begin
      mem_ctrl_amo <= ex_ctrl_amo;
    end
    if(T11) begin
      ex_ctrl_amo <= id_ctrl_amo;
    end
    if(T451) begin
      mem_ctrl_fence <= ex_ctrl_fence;
    end
    if(T11) begin
      ex_ctrl_fence <= id_ctrl_fence;
    end
    if(T451) begin
      mem_ctrl_scall <= ex_ctrl_scall;
    end
    if(T11) begin
      ex_ctrl_scall <= id_ctrl_scall;
    end
    if(T451) begin
      mem_ctrl_rfs3 <= ex_ctrl_rfs3;
    end
    if(T11) begin
      ex_ctrl_rfs3 <= id_ctrl_rfs3;
    end
    if(T451) begin
      mem_ctrl_rfs2 <= ex_ctrl_rfs2;
    end
    if(T11) begin
      ex_ctrl_rfs2 <= id_ctrl_rfs2;
    end
    if(T451) begin
      mem_ctrl_rfs1 <= ex_ctrl_rfs1;
    end
    if(T11) begin
      ex_ctrl_rfs1 <= id_ctrl_rfs1;
    end
    if(T451) begin
      mem_ctrl_mem_type <= ex_ctrl_mem_type;
    end
    if(T451) begin
      mem_ctrl_mem_cmd <= ex_ctrl_mem_cmd;
    end
    if(T451) begin
      mem_ctrl_alu_fn <= ex_ctrl_alu_fn;
    end
    if(T11) begin
      ex_ctrl_alu_fn <= id_ctrl_alu_fn;
    end
    if(T451) begin
      mem_ctrl_alu_dw <= ex_ctrl_alu_dw;
    end
    if(T11) begin
      ex_ctrl_alu_dw <= id_ctrl_alu_dw;
    end
    if(T451) begin
      mem_ctrl_sel_imm <= ex_ctrl_sel_imm;
    end
    if(T11) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if(T451) begin
      mem_ctrl_sel_alu1 <= ex_ctrl_sel_alu1;
    end
    if(T11) begin
      ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
    end
    if(T451) begin
      mem_ctrl_sel_alu2 <= ex_ctrl_sel_alu2;
    end
    if(T11) begin
      ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
    end
    if(T451) begin
      mem_ctrl_rxs1 <= ex_ctrl_rxs1;
    end
    if(T11) begin
      ex_ctrl_rxs1 <= id_ctrl_rxs1;
    end
    if(T451) begin
      mem_ctrl_rxs2 <= ex_ctrl_rxs2;
    end
    if(T11) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if(T451) begin
      mem_ctrl_legal <= ex_ctrl_legal;
    end
    if(T11) begin
      ex_ctrl_legal <= id_ctrl_legal;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T133;
  wire cmp;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] T29;
  wire T30;
  wire[63:0] shout_l;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[62:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[61:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[59:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[55:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[47:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T134;
  wire[31:0] T55;
  wire[63:0] T56;
  wire[63:0] T135;
  wire[47:0] T57;
  wire[63:0] T58;
  wire[63:0] T136;
  wire[55:0] T59;
  wire[63:0] T60;
  wire[63:0] T137;
  wire[59:0] T61;
  wire[63:0] T62;
  wire[63:0] T138;
  wire[61:0] T63;
  wire[63:0] T64;
  wire[63:0] T139;
  wire[62:0] T65;
  wire T66;
  wire[63:0] shout_r;
  wire[64:0] T67;
  wire[5:0] shamt;
  wire[5:0] T68;
  wire[4:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[64:0] T73;
  wire[64:0] T74;
  wire[63:0] shin;
  wire[63:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[62:0] T78;
  wire[63:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[61:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[59:0] T86;
  wire[63:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[55:0] T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[47:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[31:0] T98;
  wire[63:0] T99;
  wire[63:0] T140;
  wire[31:0] T100;
  wire[63:0] T101;
  wire[63:0] T141;
  wire[47:0] T102;
  wire[63:0] T103;
  wire[63:0] T142;
  wire[55:0] T104;
  wire[63:0] T105;
  wire[63:0] T143;
  wire[59:0] T106;
  wire[63:0] T107;
  wire[63:0] T144;
  wire[61:0] T108;
  wire[63:0] T109;
  wire[63:0] T145;
  wire[62:0] T110;
  wire[63:0] shin_r;
  wire[31:0] T111;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T112;
  wire[31:0] T146;
  wire T113;
  wire T114;
  wire[31:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[31:0] out_hi;
  wire[31:0] T129;
  wire[31:0] T147;
  wire T130;
  wire[31:0] T131;
  wire T132;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T126 ? sum : T6;
  assign T6 = T123 ? shout_r : T7;
  assign T7 = T66 ? shout_l : T8;
  assign T8 = T30 ? T29 : T9;
  assign T9 = T28 ? T27 : T10;
  assign T10 = T26 ? T25 : T133;
  assign T133 = {63'h0, cmp};
  assign cmp = T24 ^ T11;
  assign T11 = T22 ? T21 : T12;
  assign T12 = T18 ? T17 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = io_in1[6'h3f:6'h3f];
  assign T15 = io_in2[6'h3f:6'h3f];
  assign T16 = io_fn[1'h1:1'h1];
  assign T17 = sum[6'h3f:6'h3f];
  assign T18 = T20 == T19;
  assign T19 = io_in2[6'h3f:6'h3f];
  assign T20 = io_in1[6'h3f:6'h3f];
  assign T21 = sum == 64'h0;
  assign T22 = T23 ^ 1'h1;
  assign T23 = io_fn[2'h2:2'h2];
  assign T24 = io_fn[1'h0:1'h0];
  assign T25 = io_in1 ^ io_in2;
  assign T26 = io_fn == 4'h4;
  assign T27 = io_in1 | io_in2;
  assign T28 = io_fn == 4'h6;
  assign T29 = io_in1 & io_in2;
  assign T30 = io_fn == 4'h7;
  assign shout_l = T64 | T31;
  assign T31 = T32 & 64'haaaaaaaaaaaaaaaa;
  assign T32 = T33 << 1'h1;
  assign T33 = T34[6'h3e:1'h0];
  assign T34 = T62 | T35;
  assign T35 = T36 & 64'hcccccccccccccccc;
  assign T36 = T37 << 2'h2;
  assign T37 = T38[6'h3d:1'h0];
  assign T38 = T60 | T39;
  assign T39 = T40 & 64'hf0f0f0f0f0f0f0f0;
  assign T40 = T41 << 3'h4;
  assign T41 = T42[6'h3b:1'h0];
  assign T42 = T58 | T43;
  assign T43 = T44 & 64'hff00ff00ff00ff00;
  assign T44 = T45 << 4'h8;
  assign T45 = T46[6'h37:1'h0];
  assign T46 = T56 | T47;
  assign T47 = T48 & 64'hffff0000ffff0000;
  assign T48 = T49 << 5'h10;
  assign T49 = T50[6'h2f:1'h0];
  assign T50 = T54 | T51;
  assign T51 = T52 & 64'hffffffff00000000;
  assign T52 = T53 << 6'h20;
  assign T53 = shout_r[5'h1f:1'h0];
  assign T54 = T134 & 64'hffffffff;
  assign T134 = {32'h0, T55};
  assign T55 = shout_r >> 6'h20;
  assign T56 = T135 & 64'hffff0000ffff;
  assign T135 = {16'h0, T57};
  assign T57 = T50 >> 5'h10;
  assign T58 = T136 & 64'hff00ff00ff00ff;
  assign T136 = {8'h0, T59};
  assign T59 = T46 >> 4'h8;
  assign T60 = T137 & 64'hf0f0f0f0f0f0f0f;
  assign T137 = {4'h0, T61};
  assign T61 = T42 >> 3'h4;
  assign T62 = T138 & 64'h3333333333333333;
  assign T138 = {2'h0, T63};
  assign T63 = T38 >> 2'h2;
  assign T64 = T139 & 64'h5555555555555555;
  assign T139 = {1'h0, T65};
  assign T65 = T34 >> 1'h1;
  assign T66 = io_fn == 4'h1;
  assign shout_r = T67[6'h3f:1'h0];
  assign T67 = $signed(T73) >>> shamt;
  assign shamt = T68;
  assign T68 = {T70, T69};
  assign T69 = io_in2[3'h4:1'h0];
  assign T70 = T72 & T71;
  assign T71 = io_dw == 1'h1;
  assign T72 = io_in2[3'h5:3'h5];
  assign T73 = T74;
  assign T74 = {T120, shin};
  assign shin = T117 ? shin_r : T75;
  assign T75 = T109 | T76;
  assign T76 = T77 & 64'haaaaaaaaaaaaaaaa;
  assign T77 = T78 << 1'h1;
  assign T78 = T79[6'h3e:1'h0];
  assign T79 = T107 | T80;
  assign T80 = T81 & 64'hcccccccccccccccc;
  assign T81 = T82 << 2'h2;
  assign T82 = T83[6'h3d:1'h0];
  assign T83 = T105 | T84;
  assign T84 = T85 & 64'hf0f0f0f0f0f0f0f0;
  assign T85 = T86 << 3'h4;
  assign T86 = T87[6'h3b:1'h0];
  assign T87 = T103 | T88;
  assign T88 = T89 & 64'hff00ff00ff00ff00;
  assign T89 = T90 << 4'h8;
  assign T90 = T91[6'h37:1'h0];
  assign T91 = T101 | T92;
  assign T92 = T93 & 64'hffff0000ffff0000;
  assign T93 = T94 << 5'h10;
  assign T94 = T95[6'h2f:1'h0];
  assign T95 = T99 | T96;
  assign T96 = T97 & 64'hffffffff00000000;
  assign T97 = T98 << 6'h20;
  assign T98 = shin_r[5'h1f:1'h0];
  assign T99 = T140 & 64'hffffffff;
  assign T140 = {32'h0, T100};
  assign T100 = shin_r >> 6'h20;
  assign T101 = T141 & 64'hffff0000ffff;
  assign T141 = {16'h0, T102};
  assign T102 = T95 >> 5'h10;
  assign T103 = T142 & 64'hff00ff00ff00ff;
  assign T142 = {8'h0, T104};
  assign T104 = T91 >> 4'h8;
  assign T105 = T143 & 64'hf0f0f0f0f0f0f0f;
  assign T143 = {4'h0, T106};
  assign T106 = T87 >> 3'h4;
  assign T107 = T144 & 64'h3333333333333333;
  assign T144 = {2'h0, T108};
  assign T108 = T83 >> 2'h2;
  assign T109 = T145 & 64'h5555555555555555;
  assign T145 = {1'h0, T110};
  assign T110 = T79 >> 1'h1;
  assign shin_r = {shin_hi, T111};
  assign T111 = io_in1[5'h1f:1'h0];
  assign shin_hi = T116 ? T115 : shin_hi_32;
  assign shin_hi_32 = T114 ? T112 : 32'h0;
  assign T112 = 32'h0 - T146;
  assign T146 = {31'h0, T113};
  assign T113 = io_in1[5'h1f:5'h1f];
  assign T114 = io_fn[2'h3:2'h3];
  assign T115 = io_in1[6'h3f:6'h20];
  assign T116 = io_dw == 1'h1;
  assign T117 = T119 | T118;
  assign T118 = io_fn == 4'hb;
  assign T119 = io_fn == 4'h5;
  assign T120 = T122 & T121;
  assign T121 = shin[6'h3f:6'h3f];
  assign T122 = io_fn[2'h3:2'h3];
  assign T123 = T125 | T124;
  assign T124 = io_fn == 4'hb;
  assign T125 = io_fn == 4'h5;
  assign T126 = T128 | T127;
  assign T127 = io_fn == 4'ha;
  assign T128 = io_fn == 4'h0;
  assign out_hi = T132 ? T131 : T129;
  assign T129 = 32'h0 - T147;
  assign T147 = {31'h0, T130};
  assign T130 = out64[5'h1f:5'h1f];
  assign T131 = out64[6'h3f:6'h20];
  assign T132 = io_dw == 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[129:0] T180;
  wire[63:0] negated_remainder;
  wire[63:0] T119;
  wire T11;
  wire T12;
  reg  isMul;
  wire T13;
  wire cmdMul;
  wire T14;
  wire[3:0] T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  reg [2:0] state;
  wire[2:0] T181;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  reg  neg_out;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  isHi;
  wire T33;
  wire cmdHi;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire T37;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T41;
  wire[64:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[64:0] T46;
  wire[63:0] rhs_in;
  wire[31:0] T47;
  wire[31:0] T48;
  wire[31:0] T49;
  wire[31:0] T182;
  wire[31:0] T50;
  wire T51;
  wire rhs_sign;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire rhsSigned;
  wire T56;
  wire[3:0] T57;
  wire[64:0] T58;
  wire T59;
  reg [6:0] count;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire[6:0] T65;
  wire[6:0] T183;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[5:0] T184;
  wire[5:0] T185;
  wire[5:0] T186;
  wire[5:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[5:0] T190;
  wire[5:0] T191;
  wire[5:0] T192;
  wire[5:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire[5:0] T196;
  wire[5:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[4:0] T216;
  wire[4:0] T217;
  wire[4:0] T218;
  wire[4:0] T219;
  wire[4:0] T220;
  wire[4:0] T221;
  wire[4:0] T222;
  wire[4:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[4:0] T226;
  wire[4:0] T227;
  wire[4:0] T228;
  wire[4:0] T229;
  wire[4:0] T230;
  wire[4:0] T231;
  wire[3:0] T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[3:0] T238;
  wire[3:0] T239;
  wire[2:0] T240;
  wire[2:0] T241;
  wire[2:0] T242;
  wire[2:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire T246;
  wire[63:0] T70;
  wire[63:0] T71;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire[5:0] T72;
  wire[5:0] T309;
  wire[5:0] T310;
  wire[5:0] T311;
  wire[5:0] T312;
  wire[5:0] T313;
  wire[5:0] T314;
  wire[5:0] T315;
  wire[5:0] T316;
  wire[5:0] T317;
  wire[5:0] T318;
  wire[5:0] T319;
  wire[5:0] T320;
  wire[5:0] T321;
  wire[5:0] T322;
  wire[5:0] T323;
  wire[5:0] T324;
  wire[5:0] T325;
  wire[5:0] T326;
  wire[5:0] T327;
  wire[5:0] T328;
  wire[5:0] T329;
  wire[5:0] T330;
  wire[5:0] T331;
  wire[5:0] T332;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[4:0] T341;
  wire[4:0] T342;
  wire[4:0] T343;
  wire[4:0] T344;
  wire[4:0] T345;
  wire[4:0] T346;
  wire[4:0] T347;
  wire[4:0] T348;
  wire[4:0] T349;
  wire[4:0] T350;
  wire[4:0] T351;
  wire[4:0] T352;
  wire[4:0] T353;
  wire[4:0] T354;
  wire[4:0] T355;
  wire[4:0] T356;
  wire[3:0] T357;
  wire[3:0] T358;
  wire[3:0] T359;
  wire[3:0] T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[2:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire[2:0] T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire T371;
  wire[63:0] T74;
  wire[63:0] T75;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire lhs_sign;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire lhsSigned;
  wire T84;
  wire[3:0] T85;
  wire T86;
  wire T87;
  wire[2:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[64:0] T97;
  wire[5:0] T98;
  wire[10:0] T99;
  wire[63:0] T100;
  wire[128:0] T101;
  wire[63:0] T102;
  wire[64:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[2:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire[129:0] T434;
  wire T120;
  wire[129:0] T435;
  wire[63:0] T121;
  wire T122;
  wire[129:0] T123;
  wire[129:0] T124;
  wire[64:0] T125;
  wire[63:0] T126;
  wire[128:0] T127;
  wire[63:0] T128;
  wire[128:0] T129;
  wire[128:0] T130;
  wire[128:0] T131;
  wire[55:0] T132;
  wire[72:0] T133;
  wire[72:0] T436;
  wire[64:0] T134;
  wire[64:0] T135;
  wire[7:0] T437;
  wire T438;
  wire[72:0] T136;
  wire[8:0] T137;
  wire[8:0] T138;
  wire[7:0] T139;
  wire[64:0] T140;
  wire[128:0] T141;
  wire[5:0] T142;
  wire[10:0] T143;
  wire[10:0] T144;
  wire[64:0] T145;
  wire[64:0] T146;
  wire T147;
  wire T148;
  wire[129:0] T439;
  wire[128:0] T149;
  wire[64:0] T150;
  wire T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[63:0] T154;
  wire[63:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[129:0] T440;
  wire[126:0] T159;
  wire[63:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire[129:0] T441;
  wire[63:0] lhs_in;
  wire[31:0] T167;
  wire[31:0] T168;
  wire[31:0] T169;
  wire[31:0] T442;
  wire[31:0] T170;
  wire T171;
  wire[63:0] T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T443;
  wire T175;
  wire T176;
  reg  req_dw;
  wire T177;
  wire T178;
  wire T179;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T176 ? T172 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T441 : T5;
  assign T5 = T161 ? T440 : T6;
  assign T6 = T156 ? T439 : T7;
  assign T7 = T147 ? T123 : T8;
  assign T8 = T122 ? T435 : T9;
  assign T9 = T120 ? T434 : T10;
  assign T10 = T11 ? T180 : remainder;
  assign T180 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T119;
  assign T119 = remainder[6'h3f:1'h0];
  assign T11 = T19 & T12;
  assign T12 = T18 | isMul;
  assign T13 = T1 ? cmdMul : isMul;
  assign cmdMul = T16 | T14;
  assign T14 = T15 == 4'h8;
  assign T15 = io_req_bits_fn & 4'h8;
  assign T16 = T17 == 4'h0;
  assign T17 = io_req_bits_fn & 4'h4;
  assign T18 = remainder[6'h3f:6'h3f];
  assign T19 = state == 3'h1;
  assign T181 = reset ? 3'h0 : T20;
  assign T20 = T1 ? T115 : T21;
  assign T21 = T113 ? 3'h0 : T22;
  assign T22 = T111 ? T109 : T23;
  assign T23 = T89 ? T88 : T24;
  assign T24 = T122 ? T27 : T25;
  assign T25 = T120 ? 3'h5 : T26;
  assign T26 = T19 ? 3'h2 : state;
  assign T27 = neg_out ? 3'h4 : 3'h5;
  assign T28 = T1 ? T77 : T29;
  assign T29 = T30 ? 1'h0 : neg_out;
  assign T30 = T156 & T31;
  assign T31 = T39 & T32;
  assign T32 = isHi ^ 1'h1;
  assign T33 = T1 ? cmdHi : isHi;
  assign cmdHi = T34 | T14;
  assign T34 = T37 | T35;
  assign T35 = T36 == 4'h2;
  assign T36 = io_req_bits_fn & 4'h2;
  assign T37 = T38 == 4'h1;
  assign T38 = io_req_bits_fn & 4'h5;
  assign T39 = T59 & T40;
  assign T40 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T58 - divisor;
  assign T41 = T1 ? T46 : T42;
  assign T42 = T43 ? subtractor : divisor;
  assign T43 = T19 & T44;
  assign T44 = T45 | isMul;
  assign T45 = divisor[6'h3f:6'h3f];
  assign T46 = {rhs_sign, rhs_in};
  assign rhs_in = {T48, T47};
  assign T47 = io_req_bits_in2[5'h1f:1'h0];
  assign T48 = T51 ? T50 : T49;
  assign T49 = 32'h0 - T182;
  assign T182 = {31'h0, rhs_sign};
  assign T50 = io_req_bits_in2[6'h3f:6'h20];
  assign T51 = io_req_bits_dw == 1'h1;
  assign rhs_sign = rhsSigned & T52;
  assign T52 = T55 ? T54 : T53;
  assign T53 = io_req_bits_in2[5'h1f:5'h1f];
  assign T54 = io_req_bits_in2[6'h3f:6'h3f];
  assign T55 = io_req_bits_dw == 1'h1;
  assign rhsSigned = T56 | T16;
  assign T56 = T57 == 4'h0;
  assign T57 = io_req_bits_fn & 4'h9;
  assign T58 = remainder[8'h80:7'h40];
  assign T59 = count == 7'h0;
  assign T60 = T1 ? 7'h0 : T61;
  assign T61 = T161 ? T183 : T62;
  assign T62 = T156 ? T65 : T63;
  assign T63 = T147 ? T64 : count;
  assign T64 = count + 7'h1;
  assign T65 = count + 7'h1;
  assign T183 = {1'h0, T66};
  assign T66 = T76 ? 6'h3f : T67;
  assign T67 = T68[3'h5:1'h0];
  assign T68 = T72 - T184;
  assign T184 = T308 ? 6'h3f : T185;
  assign T185 = T307 ? 6'h3e : T186;
  assign T186 = T306 ? 6'h3d : T187;
  assign T187 = T305 ? 6'h3c : T188;
  assign T188 = T304 ? 6'h3b : T189;
  assign T189 = T303 ? 6'h3a : T190;
  assign T190 = T302 ? 6'h39 : T191;
  assign T191 = T301 ? 6'h38 : T192;
  assign T192 = T300 ? 6'h37 : T193;
  assign T193 = T299 ? 6'h36 : T194;
  assign T194 = T298 ? 6'h35 : T195;
  assign T195 = T297 ? 6'h34 : T196;
  assign T196 = T296 ? 6'h33 : T197;
  assign T197 = T295 ? 6'h32 : T198;
  assign T198 = T294 ? 6'h31 : T199;
  assign T199 = T293 ? 6'h30 : T200;
  assign T200 = T292 ? 6'h2f : T201;
  assign T201 = T291 ? 6'h2e : T202;
  assign T202 = T290 ? 6'h2d : T203;
  assign T203 = T289 ? 6'h2c : T204;
  assign T204 = T288 ? 6'h2b : T205;
  assign T205 = T287 ? 6'h2a : T206;
  assign T206 = T286 ? 6'h29 : T207;
  assign T207 = T285 ? 6'h28 : T208;
  assign T208 = T284 ? 6'h27 : T209;
  assign T209 = T283 ? 6'h26 : T210;
  assign T210 = T282 ? 6'h25 : T211;
  assign T211 = T281 ? 6'h24 : T212;
  assign T212 = T280 ? 6'h23 : T213;
  assign T213 = T279 ? 6'h22 : T214;
  assign T214 = T278 ? 6'h21 : T215;
  assign T215 = T277 ? 6'h20 : T216;
  assign T216 = T276 ? 5'h1f : T217;
  assign T217 = T275 ? 5'h1e : T218;
  assign T218 = T274 ? 5'h1d : T219;
  assign T219 = T273 ? 5'h1c : T220;
  assign T220 = T272 ? 5'h1b : T221;
  assign T221 = T271 ? 5'h1a : T222;
  assign T222 = T270 ? 5'h19 : T223;
  assign T223 = T269 ? 5'h18 : T224;
  assign T224 = T268 ? 5'h17 : T225;
  assign T225 = T267 ? 5'h16 : T226;
  assign T226 = T266 ? 5'h15 : T227;
  assign T227 = T265 ? 5'h14 : T228;
  assign T228 = T264 ? 5'h13 : T229;
  assign T229 = T263 ? 5'h12 : T230;
  assign T230 = T262 ? 5'h11 : T231;
  assign T231 = T261 ? 5'h10 : T232;
  assign T232 = T260 ? 4'hf : T233;
  assign T233 = T259 ? 4'he : T234;
  assign T234 = T258 ? 4'hd : T235;
  assign T235 = T257 ? 4'hc : T236;
  assign T236 = T256 ? 4'hb : T237;
  assign T237 = T255 ? 4'ha : T238;
  assign T238 = T254 ? 4'h9 : T239;
  assign T239 = T253 ? 4'h8 : T240;
  assign T240 = T252 ? 3'h7 : T241;
  assign T241 = T251 ? 3'h6 : T242;
  assign T242 = T250 ? 3'h5 : T243;
  assign T243 = T249 ? 3'h4 : T244;
  assign T244 = T248 ? 2'h3 : T245;
  assign T245 = T247 ? 2'h2 : T246;
  assign T246 = T70[1'h1:1'h1];
  assign T70 = T71[6'h3f:1'h0];
  assign T71 = remainder[6'h3f:1'h0];
  assign T247 = T70[2'h2:2'h2];
  assign T248 = T70[2'h3:2'h3];
  assign T249 = T70[3'h4:3'h4];
  assign T250 = T70[3'h5:3'h5];
  assign T251 = T70[3'h6:3'h6];
  assign T252 = T70[3'h7:3'h7];
  assign T253 = T70[4'h8:4'h8];
  assign T254 = T70[4'h9:4'h9];
  assign T255 = T70[4'ha:4'ha];
  assign T256 = T70[4'hb:4'hb];
  assign T257 = T70[4'hc:4'hc];
  assign T258 = T70[4'hd:4'hd];
  assign T259 = T70[4'he:4'he];
  assign T260 = T70[4'hf:4'hf];
  assign T261 = T70[5'h10:5'h10];
  assign T262 = T70[5'h11:5'h11];
  assign T263 = T70[5'h12:5'h12];
  assign T264 = T70[5'h13:5'h13];
  assign T265 = T70[5'h14:5'h14];
  assign T266 = T70[5'h15:5'h15];
  assign T267 = T70[5'h16:5'h16];
  assign T268 = T70[5'h17:5'h17];
  assign T269 = T70[5'h18:5'h18];
  assign T270 = T70[5'h19:5'h19];
  assign T271 = T70[5'h1a:5'h1a];
  assign T272 = T70[5'h1b:5'h1b];
  assign T273 = T70[5'h1c:5'h1c];
  assign T274 = T70[5'h1d:5'h1d];
  assign T275 = T70[5'h1e:5'h1e];
  assign T276 = T70[5'h1f:5'h1f];
  assign T277 = T70[6'h20:6'h20];
  assign T278 = T70[6'h21:6'h21];
  assign T279 = T70[6'h22:6'h22];
  assign T280 = T70[6'h23:6'h23];
  assign T281 = T70[6'h24:6'h24];
  assign T282 = T70[6'h25:6'h25];
  assign T283 = T70[6'h26:6'h26];
  assign T284 = T70[6'h27:6'h27];
  assign T285 = T70[6'h28:6'h28];
  assign T286 = T70[6'h29:6'h29];
  assign T287 = T70[6'h2a:6'h2a];
  assign T288 = T70[6'h2b:6'h2b];
  assign T289 = T70[6'h2c:6'h2c];
  assign T290 = T70[6'h2d:6'h2d];
  assign T291 = T70[6'h2e:6'h2e];
  assign T292 = T70[6'h2f:6'h2f];
  assign T293 = T70[6'h30:6'h30];
  assign T294 = T70[6'h31:6'h31];
  assign T295 = T70[6'h32:6'h32];
  assign T296 = T70[6'h33:6'h33];
  assign T297 = T70[6'h34:6'h34];
  assign T298 = T70[6'h35:6'h35];
  assign T299 = T70[6'h36:6'h36];
  assign T300 = T70[6'h37:6'h37];
  assign T301 = T70[6'h38:6'h38];
  assign T302 = T70[6'h39:6'h39];
  assign T303 = T70[6'h3a:6'h3a];
  assign T304 = T70[6'h3b:6'h3b];
  assign T305 = T70[6'h3c:6'h3c];
  assign T306 = T70[6'h3d:6'h3d];
  assign T307 = T70[6'h3e:6'h3e];
  assign T308 = T70[6'h3f:6'h3f];
  assign T72 = 6'h3f + T309;
  assign T309 = T433 ? 6'h3f : T310;
  assign T310 = T432 ? 6'h3e : T311;
  assign T311 = T431 ? 6'h3d : T312;
  assign T312 = T430 ? 6'h3c : T313;
  assign T313 = T429 ? 6'h3b : T314;
  assign T314 = T428 ? 6'h3a : T315;
  assign T315 = T427 ? 6'h39 : T316;
  assign T316 = T426 ? 6'h38 : T317;
  assign T317 = T425 ? 6'h37 : T318;
  assign T318 = T424 ? 6'h36 : T319;
  assign T319 = T423 ? 6'h35 : T320;
  assign T320 = T422 ? 6'h34 : T321;
  assign T321 = T421 ? 6'h33 : T322;
  assign T322 = T420 ? 6'h32 : T323;
  assign T323 = T419 ? 6'h31 : T324;
  assign T324 = T418 ? 6'h30 : T325;
  assign T325 = T417 ? 6'h2f : T326;
  assign T326 = T416 ? 6'h2e : T327;
  assign T327 = T415 ? 6'h2d : T328;
  assign T328 = T414 ? 6'h2c : T329;
  assign T329 = T413 ? 6'h2b : T330;
  assign T330 = T412 ? 6'h2a : T331;
  assign T331 = T411 ? 6'h29 : T332;
  assign T332 = T410 ? 6'h28 : T333;
  assign T333 = T409 ? 6'h27 : T334;
  assign T334 = T408 ? 6'h26 : T335;
  assign T335 = T407 ? 6'h25 : T336;
  assign T336 = T406 ? 6'h24 : T337;
  assign T337 = T405 ? 6'h23 : T338;
  assign T338 = T404 ? 6'h22 : T339;
  assign T339 = T403 ? 6'h21 : T340;
  assign T340 = T402 ? 6'h20 : T341;
  assign T341 = T401 ? 5'h1f : T342;
  assign T342 = T400 ? 5'h1e : T343;
  assign T343 = T399 ? 5'h1d : T344;
  assign T344 = T398 ? 5'h1c : T345;
  assign T345 = T397 ? 5'h1b : T346;
  assign T346 = T396 ? 5'h1a : T347;
  assign T347 = T395 ? 5'h19 : T348;
  assign T348 = T394 ? 5'h18 : T349;
  assign T349 = T393 ? 5'h17 : T350;
  assign T350 = T392 ? 5'h16 : T351;
  assign T351 = T391 ? 5'h15 : T352;
  assign T352 = T390 ? 5'h14 : T353;
  assign T353 = T389 ? 5'h13 : T354;
  assign T354 = T388 ? 5'h12 : T355;
  assign T355 = T387 ? 5'h11 : T356;
  assign T356 = T386 ? 5'h10 : T357;
  assign T357 = T385 ? 4'hf : T358;
  assign T358 = T384 ? 4'he : T359;
  assign T359 = T383 ? 4'hd : T360;
  assign T360 = T382 ? 4'hc : T361;
  assign T361 = T381 ? 4'hb : T362;
  assign T362 = T380 ? 4'ha : T363;
  assign T363 = T379 ? 4'h9 : T364;
  assign T364 = T378 ? 4'h8 : T365;
  assign T365 = T377 ? 3'h7 : T366;
  assign T366 = T376 ? 3'h6 : T367;
  assign T367 = T375 ? 3'h5 : T368;
  assign T368 = T374 ? 3'h4 : T369;
  assign T369 = T373 ? 2'h3 : T370;
  assign T370 = T372 ? 2'h2 : T371;
  assign T371 = T74[1'h1:1'h1];
  assign T74 = T75[6'h3f:1'h0];
  assign T75 = divisor[6'h3f:1'h0];
  assign T372 = T74[2'h2:2'h2];
  assign T373 = T74[2'h3:2'h3];
  assign T374 = T74[3'h4:3'h4];
  assign T375 = T74[3'h5:3'h5];
  assign T376 = T74[3'h6:3'h6];
  assign T377 = T74[3'h7:3'h7];
  assign T378 = T74[4'h8:4'h8];
  assign T379 = T74[4'h9:4'h9];
  assign T380 = T74[4'ha:4'ha];
  assign T381 = T74[4'hb:4'hb];
  assign T382 = T74[4'hc:4'hc];
  assign T383 = T74[4'hd:4'hd];
  assign T384 = T74[4'he:4'he];
  assign T385 = T74[4'hf:4'hf];
  assign T386 = T74[5'h10:5'h10];
  assign T387 = T74[5'h11:5'h11];
  assign T388 = T74[5'h12:5'h12];
  assign T389 = T74[5'h13:5'h13];
  assign T390 = T74[5'h14:5'h14];
  assign T391 = T74[5'h15:5'h15];
  assign T392 = T74[5'h16:5'h16];
  assign T393 = T74[5'h17:5'h17];
  assign T394 = T74[5'h18:5'h18];
  assign T395 = T74[5'h19:5'h19];
  assign T396 = T74[5'h1a:5'h1a];
  assign T397 = T74[5'h1b:5'h1b];
  assign T398 = T74[5'h1c:5'h1c];
  assign T399 = T74[5'h1d:5'h1d];
  assign T400 = T74[5'h1e:5'h1e];
  assign T401 = T74[5'h1f:5'h1f];
  assign T402 = T74[6'h20:6'h20];
  assign T403 = T74[6'h21:6'h21];
  assign T404 = T74[6'h22:6'h22];
  assign T405 = T74[6'h23:6'h23];
  assign T406 = T74[6'h24:6'h24];
  assign T407 = T74[6'h25:6'h25];
  assign T408 = T74[6'h26:6'h26];
  assign T409 = T74[6'h27:6'h27];
  assign T410 = T74[6'h28:6'h28];
  assign T411 = T74[6'h29:6'h29];
  assign T412 = T74[6'h2a:6'h2a];
  assign T413 = T74[6'h2b:6'h2b];
  assign T414 = T74[6'h2c:6'h2c];
  assign T415 = T74[6'h2d:6'h2d];
  assign T416 = T74[6'h2e:6'h2e];
  assign T417 = T74[6'h2f:6'h2f];
  assign T418 = T74[6'h30:6'h30];
  assign T419 = T74[6'h31:6'h31];
  assign T420 = T74[6'h32:6'h32];
  assign T421 = T74[6'h33:6'h33];
  assign T422 = T74[6'h34:6'h34];
  assign T423 = T74[6'h35:6'h35];
  assign T424 = T74[6'h36:6'h36];
  assign T425 = T74[6'h37:6'h37];
  assign T426 = T74[6'h38:6'h38];
  assign T427 = T74[6'h39:6'h39];
  assign T428 = T74[6'h3a:6'h3a];
  assign T429 = T74[6'h3b:6'h3b];
  assign T430 = T74[6'h3c:6'h3c];
  assign T431 = T74[6'h3d:6'h3d];
  assign T432 = T74[6'h3e:6'h3e];
  assign T433 = T74[6'h3f:6'h3f];
  assign T76 = T184 < T309;
  assign T77 = T87 & T78;
  assign T78 = cmdHi ? lhs_sign : T79;
  assign T79 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T80;
  assign T80 = T83 ? T82 : T81;
  assign T81 = io_req_bits_in1[5'h1f:5'h1f];
  assign T82 = io_req_bits_in1[6'h3f:6'h3f];
  assign T83 = io_req_bits_dw == 1'h1;
  assign lhsSigned = T86 | T84;
  assign T84 = T85 == 4'h0;
  assign T85 = io_req_bits_fn & 4'h3;
  assign T86 = T56 | T16;
  assign T87 = cmdMul ^ 1'h1;
  assign T88 = isHi ? 3'h3 : 3'h5;
  assign T89 = T147 & T90;
  assign T90 = T92 | T91;
  assign T91 = count == 7'h7;
  assign T92 = T104 & T93;
  assign T93 = T94 == 64'h0;
  assign T94 = T100 & T95;
  assign T95 = ~ T96;
  assign T96 = T97[6'h3f:1'h0];
  assign T97 = $signed(65'h10000000000000000) >>> T98;
  assign T98 = T99[3'h5:1'h0];
  assign T99 = count * 4'h8;
  assign T100 = T101[6'h3f:1'h0];
  assign T101 = {T103, T102};
  assign T102 = remainder[6'h3f:1'h0];
  assign T103 = remainder[8'h81:7'h41];
  assign T104 = T106 & T105;
  assign T105 = isHi ^ 1'h1;
  assign T106 = T108 & T107;
  assign T107 = count != 7'h0;
  assign T108 = count != 7'h7;
  assign T109 = isHi ? 3'h3 : T110;
  assign T110 = neg_out ? 3'h4 : 3'h5;
  assign T111 = T156 & T112;
  assign T112 = count == 7'h40;
  assign T113 = T114 | io_kill;
  assign T114 = io_resp_ready & io_resp_valid;
  assign T115 = T116 ? 3'h1 : 3'h2;
  assign T116 = lhs_sign | T117;
  assign T117 = rhs_sign & T118;
  assign T118 = cmdMul ^ 1'h1;
  assign T434 = {66'h0, negated_remainder};
  assign T120 = state == 3'h4;
  assign T435 = {66'h0, T121};
  assign T121 = remainder[8'h80:7'h41];
  assign T122 = state == 3'h3;
  assign T123 = T124;
  assign T124 = {T146, T125};
  assign T125 = {1'h0, T126};
  assign T126 = T127[6'h3f:1'h0];
  assign T127 = {T145, T128};
  assign T128 = T129[6'h3f:1'h0];
  assign T129 = T92 ? T141 : T130;
  assign T130 = T131;
  assign T131 = {T133, T132};
  assign T132 = T100[6'h3f:4'h8];
  assign T133 = T136 + T436;
  assign T436 = {T437, T134};
  assign T134 = T135;
  assign T135 = T101[8'h80:7'h40];
  assign T437 = T438 ? 8'hff : 8'h0;
  assign T438 = T134[7'h40:7'h40];
  assign T136 = $signed(T140) * $signed(T137);
  assign T137 = T138;
  assign T138 = {1'h0, T139};
  assign T139 = T100[3'h7:1'h0];
  assign T140 = divisor;
  assign T141 = T101 >> T142;
  assign T142 = T143[3'h5:1'h0];
  assign T143 = 11'h40 - T144;
  assign T144 = count * 4'h8;
  assign T145 = T130[8'h80:7'h40];
  assign T146 = T127 >> 7'h40;
  assign T147 = T148 & isMul;
  assign T148 = state == 3'h2;
  assign T439 = {1'h0, T149};
  assign T149 = {T153, T150};
  assign T150 = {T152, T151};
  assign T151 = less ^ 1'h1;
  assign T152 = remainder[6'h3f:1'h0];
  assign T153 = less ? T155 : T154;
  assign T154 = subtractor[6'h3f:1'h0];
  assign T155 = remainder[7'h7f:7'h40];
  assign T156 = T158 & T157;
  assign T157 = isMul ^ 1'h1;
  assign T158 = state == 3'h2;
  assign T440 = {3'h0, T159};
  assign T159 = T160 << T66;
  assign T160 = remainder[6'h3f:1'h0];
  assign T161 = T156 & T162;
  assign T162 = T165 & T163;
  assign T163 = T164 | T76;
  assign T164 = 6'h0 < T68;
  assign T165 = T166 & less;
  assign T166 = count == 7'h0;
  assign T441 = {66'h0, lhs_in};
  assign lhs_in = {T168, T167};
  assign T167 = io_req_bits_in1[5'h1f:1'h0];
  assign T168 = T171 ? T170 : T169;
  assign T169 = 32'h0 - T442;
  assign T442 = {31'h0, lhs_sign};
  assign T170 = io_req_bits_in1[6'h3f:6'h20];
  assign T171 = io_req_bits_dw == 1'h1;
  assign T172 = {T174, T173};
  assign T173 = remainder[5'h1f:1'h0];
  assign T174 = 32'h0 - T443;
  assign T443 = {31'h0, T175};
  assign T175 = remainder[5'h1f:5'h1f];
  assign T176 = req_dw == 1'h0;
  assign T177 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T178;
  assign T178 = state == 3'h5;
  assign io_req_ready = T179;
  assign T179 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T441;
    end else if(T161) begin
      remainder <= T440;
    end else if(T156) begin
      remainder <= T439;
    end else if(T147) begin
      remainder <= T123;
    end else if(T122) begin
      remainder <= T435;
    end else if(T120) begin
      remainder <= T434;
    end else if(T11) begin
      remainder <= T180;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T115;
    end else if(T113) begin
      state <= 3'h0;
    end else if(T111) begin
      state <= T109;
    end else if(T89) begin
      state <= T88;
    end else if(T122) begin
      state <= T27;
    end else if(T120) begin
      state <= 3'h5;
    end else if(T19) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T77;
    end else if(T30) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T46;
    end else if(T43) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T161) begin
      count <= T183;
    end else if(T156) begin
      count <= T65;
    end else if(T147) begin
      count <= T64;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [1:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output[7:0] io_status_ip,
    output[7:0] io_status_im,
    output[6:0] io_status_zero,
    output io_status_er,
    output io_status_vm,
    output io_status_s64,
    output io_status_u64,
    output io_status_ef,
    output io_status_pei,
    output io_status_ei,
    output io_status_ps,
    output io_status_s,
    output[31:0] io_ptbr,
    output[43:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input  io_badvaddr_wen,
    input [43:0] io_pc,
    input  io_sret,
    output io_fatc,
    output io_replay,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [3:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[3:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[135:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_manager_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_manager_xact_id,
    //output io_rocc_dmem_acquire_ready
    input  io_rocc_dmem_acquire_valid,
    input [1:0] io_rocc_dmem_acquire_bits_header_src,
    input [1:0] io_rocc_dmem_acquire_bits_header_dst,
    input [25:0] io_rocc_dmem_acquire_bits_payload_addr,
    input [1:0] io_rocc_dmem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_acquire_bits_payload_data,
    input  io_rocc_dmem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_dmem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_dmem_acquire_bits_payload_subblock,
    input  io_rocc_dmem_grant_ready,
    //output io_rocc_dmem_grant_valid
    //output[1:0] io_rocc_dmem_grant_bits_header_src
    //output[1:0] io_rocc_dmem_grant_bits_header_dst
    //output[135:0] io_rocc_dmem_grant_bits_payload_data
    //output[1:0] io_rocc_dmem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_dmem_grant_bits_payload_manager_xact_id
    //output io_rocc_dmem_grant_bits_payload_uncached
    //output[1:0] io_rocc_dmem_grant_bits_payload_g_type
    //output io_rocc_dmem_finish_ready
    input  io_rocc_dmem_finish_valid,
    input [1:0] io_rocc_dmem_finish_bits_header_src,
    input [1:0] io_rocc_dmem_finish_bits_header_dst,
    input [3:0] io_rocc_dmem_finish_bits_payload_manager_xact_id,
    input  io_rocc_dmem_probe_ready,
    //output io_rocc_dmem_probe_valid
    //output[1:0] io_rocc_dmem_probe_bits_header_src
    //output[1:0] io_rocc_dmem_probe_bits_header_dst
    //output[25:0] io_rocc_dmem_probe_bits_payload_addr
    //output[1:0] io_rocc_dmem_probe_bits_payload_p_type
    //output io_rocc_dmem_release_ready
    input  io_rocc_dmem_release_valid,
    input [1:0] io_rocc_dmem_release_bits_header_src,
    input [1:0] io_rocc_dmem_release_bits_header_dst,
    input [25:0] io_rocc_dmem_release_bits_payload_addr,
    input [1:0] io_rocc_dmem_release_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_release_bits_payload_data,
    input [2:0] io_rocc_dmem_release_bits_payload_r_type,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  reg [2:0] reg_frm;
  wire[2:0] T479;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T480;
  wire[63:0] wdata;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T2;
  wire[63:0] T3;
  wire T4;
  wire host_pcr_req_fire;
  wire T5;
  reg  host_pcr_req_valid;
  wire T6;
  wire T7;
  wire cpu_req_valid;
  wire T8;
  wire T9;
  reg [42:0] T10;
  wire[11:0] addr;
  wire[11:0] T481;
  wire[10:0] T12;
  wire[10:0] T482;
  reg [4:0] host_pcr_bits_addr;
  wire[4:0] T13;
  wire wen;
  wire T14;
  reg  host_pcr_bits_rw;
  wire T15;
  wire[63:0] T483;
  wire[58:0] T16;
  wire T17;
  wire T18;
  wire[63:0] T19;
  reg [5:0] R20;
  wire[5:0] T484;
  wire[5:0] T21;
  wire[5:0] T22;
  wire[6:0] T23;
  wire[6:0] T485;
  wire[5:0] T24;
  wire[63:0] T25;
  wire T26;
  wire T27;
  reg [57:0] R28;
  wire[57:0] T486;
  wire[57:0] T29;
  wire[57:0] T30;
  wire[57:0] T31;
  wire T32;
  wire[57:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[43:0] T38;
  wire[43:0] T39;
  reg [43:0] reg_epc;
  wire[43:0] T40;
  wire[43:0] T41;
  wire[43:0] T42;
  wire[43:0] T43;
  wire[43:0] T44;
  wire T45;
  wire T46;
  wire[43:0] T487;
  wire[42:0] T47;
  reg [42:0] reg_evec;
  wire[42:0] T48;
  wire[42:0] T49;
  wire[42:0] T50;
  wire T51;
  wire T52;
  wire T488;
  reg [31:0] reg_ptbr;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[18:0] T56;
  wire T57;
  wire T58;
  reg  reg_status_s;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  reg_status_ps;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg  reg_status_ei;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  reg_status_pei;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg  reg_status_ef;
  wire T79;
  wire T80;
  wire T81;
  reg  reg_status_u64;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  reg  reg_status_s64;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  reg_status_vm;
  wire T90;
  wire T91;
  wire T92;
  reg  reg_status_er;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  reg [6:0] reg_status_zero;
  wire[6:0] T97;
  wire[6:0] T98;
  wire[6:0] T99;
  wire[6:0] T100;
  reg [7:0] reg_status_im;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[3:0] T105;
  wire[1:0] T106;
  reg  r_irq_ipi;
  wire T489;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[1:0] T112;
  wire T113;
  reg [63:0] reg_fromhost;
  wire[63:0] T490;
  wire[63:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg  r_irq_timer;
  wire T491;
  wire T121;
  wire T122;
  wire T123;
  reg [31:0] reg_compare;
  wire[31:0] T124;
  wire[31:0] T125;
  wire[31:0] T126;
  wire[31:0] T127;
  wire T128;
  wire T129;
  wire[63:0] T130;
  wire[63:0] T131;
  wire[63:0] T132;
  reg [5:0] R133;
  wire[5:0] T492;
  wire[5:0] T134;
  wire[5:0] T135;
  wire[6:0] T136;
  wire[6:0] T493;
  wire T137;
  reg [57:0] R138;
  wire[57:0] T494;
  wire[57:0] T139;
  wire[57:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[63:0] T144;
  wire[63:0] T145;
  wire[63:0] T146;
  reg [5:0] R147;
  wire[5:0] T495;
  wire[5:0] T148;
  wire[5:0] T149;
  wire[6:0] T150;
  wire[6:0] T496;
  wire T151;
  reg [57:0] R152;
  wire[57:0] T497;
  wire[57:0] T153;
  wire[57:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire[63:0] T158;
  wire[63:0] T159;
  wire[63:0] T160;
  reg [5:0] R161;
  wire[5:0] T498;
  wire[5:0] T162;
  wire[5:0] T163;
  wire[6:0] T164;
  wire[6:0] T499;
  wire T165;
  reg [57:0] R166;
  wire[57:0] T500;
  wire[57:0] T167;
  wire[57:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[63:0] T174;
  reg [5:0] R175;
  wire[5:0] T501;
  wire[5:0] T176;
  wire[5:0] T177;
  wire[6:0] T178;
  wire[6:0] T502;
  wire T179;
  reg [57:0] R180;
  wire[57:0] T503;
  wire[57:0] T181;
  wire[57:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire[63:0] T186;
  wire[63:0] T187;
  wire[63:0] T188;
  reg [5:0] R189;
  wire[5:0] T504;
  wire[5:0] T190;
  wire[5:0] T191;
  wire[6:0] T192;
  wire[6:0] T505;
  wire T193;
  reg [57:0] R194;
  wire[57:0] T506;
  wire[57:0] T195;
  wire[57:0] T196;
  wire T197;
  wire T198;
  wire T199;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  reg [5:0] R203;
  wire[5:0] T507;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[6:0] T206;
  wire[6:0] T508;
  wire T207;
  reg [57:0] R208;
  wire[57:0] T509;
  wire[57:0] T209;
  wire[57:0] T210;
  wire T211;
  wire T212;
  wire T213;
  wire[63:0] T214;
  wire[63:0] T215;
  wire[63:0] T216;
  reg [5:0] R217;
  wire[5:0] T510;
  wire[5:0] T218;
  wire[5:0] T219;
  wire[6:0] T220;
  wire[6:0] T511;
  wire T221;
  reg [57:0] R222;
  wire[57:0] T512;
  wire[57:0] T223;
  wire[57:0] T224;
  wire T225;
  wire T226;
  wire T227;
  wire[63:0] T228;
  wire[63:0] T229;
  wire[63:0] T230;
  reg [5:0] R231;
  wire[5:0] T513;
  wire[5:0] T232;
  wire[5:0] T233;
  wire[6:0] T234;
  wire[6:0] T514;
  wire T235;
  reg [57:0] R236;
  wire[57:0] T515;
  wire[57:0] T237;
  wire[57:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire[63:0] T242;
  wire[63:0] T243;
  wire[63:0] T244;
  reg [5:0] R245;
  wire[5:0] T516;
  wire[5:0] T246;
  wire[5:0] T247;
  wire[6:0] T248;
  wire[6:0] T517;
  wire T249;
  reg [57:0] R250;
  wire[57:0] T518;
  wire[57:0] T251;
  wire[57:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire[63:0] T256;
  wire[63:0] T257;
  wire[63:0] T258;
  reg [5:0] R259;
  wire[5:0] T519;
  wire[5:0] T260;
  wire[5:0] T261;
  wire[6:0] T262;
  wire[6:0] T520;
  wire T263;
  reg [57:0] R264;
  wire[57:0] T521;
  wire[57:0] T265;
  wire[57:0] T266;
  wire T267;
  wire T268;
  wire T269;
  wire[63:0] T270;
  wire[63:0] T271;
  wire[63:0] T272;
  reg [5:0] R273;
  wire[5:0] T522;
  wire[5:0] T274;
  wire[5:0] T275;
  wire[6:0] T276;
  wire[6:0] T523;
  wire T277;
  reg [57:0] R278;
  wire[57:0] T524;
  wire[57:0] T279;
  wire[57:0] T280;
  wire T281;
  wire T282;
  wire T283;
  wire[63:0] T284;
  wire[63:0] T285;
  wire[63:0] T286;
  reg [5:0] R287;
  wire[5:0] T525;
  wire[5:0] T288;
  wire[5:0] T289;
  wire[6:0] T290;
  wire[6:0] T526;
  wire T291;
  reg [57:0] R292;
  wire[57:0] T527;
  wire[57:0] T293;
  wire[57:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire[63:0] T298;
  wire[63:0] T299;
  wire[63:0] T300;
  reg [5:0] R301;
  wire[5:0] T528;
  wire[5:0] T302;
  wire[5:0] T303;
  wire[6:0] T304;
  wire[6:0] T529;
  wire T305;
  reg [57:0] R306;
  wire[57:0] T530;
  wire[57:0] T307;
  wire[57:0] T308;
  wire T309;
  wire T310;
  wire T311;
  wire[63:0] T312;
  wire[63:0] T313;
  wire[63:0] T314;
  reg [5:0] R315;
  wire[5:0] T531;
  wire[5:0] T316;
  wire[5:0] T317;
  wire[6:0] T318;
  wire[6:0] T532;
  wire T319;
  reg [57:0] R320;
  wire[57:0] T533;
  wire[57:0] T321;
  wire[57:0] T322;
  wire T323;
  wire T324;
  wire T325;
  wire[63:0] T326;
  wire[63:0] T327;
  wire[63:0] T328;
  reg [5:0] R329;
  wire[5:0] T534;
  wire[5:0] T330;
  wire[5:0] T331;
  wire[6:0] T332;
  wire[6:0] T535;
  wire T333;
  reg [57:0] R334;
  wire[57:0] T536;
  wire[57:0] T335;
  wire[57:0] T336;
  wire T337;
  wire T338;
  wire T339;
  wire[63:0] T340;
  wire[63:0] T341;
  wire[63:0] T342;
  reg [5:0] R343;
  wire[5:0] T537;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[6:0] T346;
  wire[6:0] T538;
  wire T347;
  reg [57:0] R348;
  wire[57:0] T539;
  wire[57:0] T349;
  wire[57:0] T350;
  wire T351;
  wire T352;
  wire T353;
  wire[63:0] T354;
  wire[63:0] T355;
  wire[63:0] T356;
  wire[63:0] T357;
  reg [63:0] reg_tohost;
  wire[63:0] T540;
  wire[63:0] T358;
  wire[63:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[63:0] T368;
  wire[63:0] T541;
  wire T369;
  reg  reg_stats;
  wire T542;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire[63:0] T374;
  wire[63:0] T543;
  wire[1:0] T375;
  wire[63:0] T376;
  wire[63:0] T544;
  wire[1:0] T377;
  wire T378;
  wire[63:0] T379;
  wire[63:0] T545;
  wire[1:0] T380;
  wire[63:0] T381;
  wire[63:0] T546;
  wire[1:0] T382;
  wire T383;
  wire[63:0] T384;
  wire[63:0] T547;
  wire T385;
  wire T386;
  wire[63:0] T387;
  wire[63:0] T548;
  wire[31:0] T388;
  wire[31:0] T389;
  wire[31:0] T390;
  wire[5:0] T391;
  wire[2:0] T392;
  wire[1:0] T393;
  wire[2:0] T394;
  wire[1:0] T395;
  wire[25:0] T396;
  wire[2:0] T397;
  wire[1:0] T398;
  wire[22:0] T399;
  wire[14:0] T400;
  wire[63:0] T401;
  wire[63:0] T402;
  reg [63:0] reg_cause;
  wire[63:0] T403;
  wire T404;
  wire[63:0] T405;
  wire[63:0] T549;
  wire[42:0] T406;
  wire[63:0] T407;
  wire[63:0] T550;
  wire[31:0] T408;
  wire[63:0] T409;
  wire[63:0] T410;
  wire[63:0] T411;
  wire[63:0] T412;
  wire[63:0] T551;
  wire[31:0] T413;
  wire[31:0] read_ptbr;
  wire[18:0] T414;
  wire[63:0] T415;
  wire[63:0] T552;
  wire[42:0] T416;
  reg [42:0] reg_badvaddr;
  wire[42:0] T553;
  wire[43:0] T417;
  wire[43:0] T554;
  wire[43:0] T418;
  wire[43:0] T419;
  wire[42:0] T420;
  wire T421;
  wire T422;
  wire[20:0] T423;
  wire T424;
  wire T425;
  wire[42:0] T426;
  wire T427;
  wire[63:0] T428;
  wire[63:0] T555;
  wire[43:0] T429;
  wire[63:0] T430;
  wire[63:0] T431;
  reg [63:0] reg_sup1;
  wire[63:0] T432;
  wire T433;
  wire T434;
  wire[63:0] T435;
  wire[63:0] T436;
  reg [63:0] reg_sup0;
  wire[63:0] T437;
  wire T438;
  wire T439;
  wire[63:0] T440;
  wire[63:0] T441;
  wire[63:0] T442;
  reg [5:0] R443;
  wire[5:0] T556;
  wire[5:0] T444;
  wire[5:0] T445;
  wire[6:0] T446;
  wire[6:0] T557;
  wire T447;
  reg [57:0] R448;
  wire[57:0] T558;
  wire[57:0] T449;
  wire[57:0] T450;
  wire T451;
  wire T452;
  wire T453;
  wire[63:0] T454;
  wire[63:0] T455;
  wire T456;
  wire[63:0] T457;
  wire[63:0] T458;
  wire T459;
  wire[63:0] T559;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  reg [4:0] reg_fflags;
  wire[4:0] T560;
  wire[63:0] T463;
  wire[63:0] T464;
  wire[63:0] T561;
  wire[4:0] T465;
  wire[4:0] T466;
  wire T467;
  wire T468;
  wire[7:0] T562;
  wire[4:0] T469;
  wire[4:0] T563;
  wire[2:0] T470;
  wire[4:0] T471;
  wire T564;
  wire T472;
  reg  host_pcr_rep_valid;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    reg_frm = {1{$random}};
    host_pcr_bits_data = {2{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    R20 = {1{$random}};
    R28 = {2{$random}};
    reg_epc = {2{$random}};
    reg_evec = {2{$random}};
    reg_ptbr = {1{$random}};
    reg_status_s = {1{$random}};
    reg_status_ps = {1{$random}};
    reg_status_ei = {1{$random}};
    reg_status_pei = {1{$random}};
    reg_status_ef = {1{$random}};
    reg_status_u64 = {1{$random}};
    reg_status_s64 = {1{$random}};
    reg_status_vm = {1{$random}};
    reg_status_er = {1{$random}};
    reg_status_zero = {1{$random}};
    reg_status_im = {1{$random}};
    r_irq_ipi = {1{$random}};
    reg_fromhost = {2{$random}};
    r_irq_timer = {1{$random}};
    reg_compare = {1{$random}};
    R133 = {1{$random}};
    R138 = {2{$random}};
    R147 = {1{$random}};
    R152 = {2{$random}};
    R161 = {1{$random}};
    R166 = {2{$random}};
    R175 = {1{$random}};
    R180 = {2{$random}};
    R189 = {1{$random}};
    R194 = {2{$random}};
    R203 = {1{$random}};
    R208 = {2{$random}};
    R217 = {1{$random}};
    R222 = {2{$random}};
    R231 = {1{$random}};
    R236 = {2{$random}};
    R245 = {1{$random}};
    R250 = {2{$random}};
    R259 = {1{$random}};
    R264 = {2{$random}};
    R273 = {1{$random}};
    R278 = {2{$random}};
    R287 = {1{$random}};
    R292 = {2{$random}};
    R301 = {1{$random}};
    R306 = {2{$random}};
    R315 = {1{$random}};
    R320 = {2{$random}};
    R329 = {1{$random}};
    R334 = {2{$random}};
    R343 = {1{$random}};
    R348 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_cause = {2{$random}};
    reg_badvaddr = {2{$random}};
    reg_sup1 = {2{$random}};
    reg_sup0 = {2{$random}};
    R443 = {1{$random}};
    R448 = {2{$random}};
    reg_fflags = {1{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
// synthesis translate_on
`endif

//  assign io_rocc_exception = {1{$random}};
//  assign io_rocc_pptw_sret = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_s = {1{$random}};
//  assign io_rocc_pptw_status_ps = {1{$random}};
//  assign io_rocc_pptw_status_ei = {1{$random}};
//  assign io_rocc_pptw_status_pei = {1{$random}};
//  assign io_rocc_pptw_status_ef = {1{$random}};
//  assign io_rocc_pptw_status_u64 = {1{$random}};
//  assign io_rocc_pptw_status_s64 = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_er = {1{$random}};
//  assign io_rocc_pptw_status_zero = {1{$random}};
//  assign io_rocc_pptw_status_im = {1{$random}};
//  assign io_rocc_pptw_status_ip = {1{$random}};
//  assign io_rocc_pptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_pptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_sret = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_s = {1{$random}};
//  assign io_rocc_dptw_status_ps = {1{$random}};
//  assign io_rocc_dptw_status_ei = {1{$random}};
//  assign io_rocc_dptw_status_pei = {1{$random}};
//  assign io_rocc_dptw_status_ef = {1{$random}};
//  assign io_rocc_dptw_status_u64 = {1{$random}};
//  assign io_rocc_dptw_status_s64 = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_er = {1{$random}};
//  assign io_rocc_dptw_status_zero = {1{$random}};
//  assign io_rocc_dptw_status_im = {1{$random}};
//  assign io_rocc_dptw_status_ip = {1{$random}};
//  assign io_rocc_dptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_dptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_sret = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_s = {1{$random}};
//  assign io_rocc_iptw_status_ps = {1{$random}};
//  assign io_rocc_iptw_status_ei = {1{$random}};
//  assign io_rocc_iptw_status_pei = {1{$random}};
//  assign io_rocc_iptw_status_ef = {1{$random}};
//  assign io_rocc_iptw_status_u64 = {1{$random}};
//  assign io_rocc_iptw_status_s64 = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_er = {1{$random}};
//  assign io_rocc_iptw_status_zero = {1{$random}};
//  assign io_rocc_iptw_status_im = {1{$random}};
//  assign io_rocc_iptw_status_ip = {1{$random}};
//  assign io_rocc_iptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_iptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_release_ready = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_p_type = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_addr = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_probe_valid = {1{$random}};
//  assign io_rocc_dmem_finish_ready = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_dmem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_grant_valid = {1{$random}};
//  assign io_rocc_dmem_acquire_ready = {1{$random}};
//  assign io_rocc_imem_finish_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_imem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_imem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
//  assign io_rocc_s = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_ptw_req_bits = {1{$random}};
//  assign io_rocc_mem_ptw_req_valid = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_data_subword = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_rocc_cmd_bits_rs2 = {2{$random}};
//  assign io_rocc_cmd_bits_rs1 = {2{$random}};
//  assign io_rocc_cmd_bits_inst_opcode = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_funct = {1{$random}};
//  assign io_rocc_cmd_valid = {1{$random}};
  assign io_fcsr_rm = reg_frm;
  assign T479 = T0[2'h2:1'h0];
  assign T0 = T17 ? T483 : T1;
  assign T1 = T8 ? wdata : T480;
  assign T480 = {61'h0, reg_frm};
  assign wdata = cpu_req_valid ? io_rw_wdata : host_pcr_bits_data;
  assign T2 = host_pcr_req_fire ? io_rw_rdata : T3;
  assign T3 = T4 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T4 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign host_pcr_req_fire = host_pcr_req_valid & T5;
  assign T5 = cpu_req_valid ^ 1'h1;
  assign T6 = host_pcr_req_fire ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : host_pcr_req_valid;
  assign cpu_req_valid = io_rw_cmd != 2'h0;
  assign T8 = wen & T9;
  assign T9 = T10[1'h1:1'h1];
  always @(*) case (addr)
    1: T10 = 43'h1;
    2: T10 = 43'h2;
    3: T10 = 43'h4;
    192: T10 = 43'h8;
    1280: T10 = 43'h10;
    1281: T10 = 43'h20;
    1282: T10 = 43'h40;
    1283: T10 = 43'h80;
    1284: T10 = 43'h100;
    1285: T10 = 43'h200;
    1286: T10 = 43'h400;
    1287: T10 = 43'h800;
    1288: T10 = 43'h1000;
    1289: T10 = 43'h2000;
    1290: T10 = 43'h4000;
    1291: T10 = 43'h8000;
    1292: T10 = 43'h10000;
    1293: T10 = 43'h20000;
    1294: T10 = 43'h40000;
    1295: T10 = 43'h80000;
    1309: T10 = 43'h100000;
    1310: T10 = 43'h200000;
    1311: T10 = 43'h400000;
    1312: T10 = 43'h800000;
    3072: T10 = 43'h1000000;
    3073: T10 = 43'h2000000;
    3074: T10 = 43'h4000000;
    3264: T10 = 43'h8000000;
    3265: T10 = 43'h10000000;
    3266: T10 = 43'h20000000;
    3267: T10 = 43'h40000000;
    3268: T10 = 43'h80000000;
    3269: T10 = 43'h100000000;
    3270: T10 = 43'h200000000;
    3271: T10 = 43'h400000000;
    3272: T10 = 43'h800000000;
    3273: T10 = 43'h1000000000;
    3274: T10 = 43'h2000000000;
    3275: T10 = 43'h4000000000;
    3276: T10 = 43'h8000000000;
    3277: T10 = 43'h10000000000;
    3278: T10 = 43'h20000000000;
    3279: T10 = 43'h40000000000;
    default: begin
      T10 = 43'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T10 = {2{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign addr = cpu_req_valid ? io_rw_addr : T481;
  assign T481 = {1'h0, T12};
  assign T12 = T482 | 11'h500;
  assign T482 = {6'h0, host_pcr_bits_addr};
  assign T13 = T4 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign wen = cpu_req_valid | T14;
  assign T14 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T15 = T4 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign T483 = {5'h0, T16};
  assign T16 = wdata >> 3'h5;
  assign T17 = wen & T18;
  assign T18 = T10[2'h2:2'h2];
  assign io_time = T19;
  assign T19 = {R28, R20};
  assign T484 = reset ? 6'h0 : T21;
  assign T21 = T26 ? T24 : T22;
  assign T22 = T23[3'h5:1'h0];
  assign T23 = T485 + 7'h1;
  assign T485 = {1'h0, R20};
  assign T24 = T25[3'h5:1'h0];
  assign T25 = wdata;
  assign T26 = wen & T27;
  assign T27 = T10[4'ha:4'ha];
  assign T486 = reset ? 58'h0 : T29;
  assign T29 = T26 ? T33 : T30;
  assign T30 = T32 ? T31 : R28;
  assign T31 = R28 + 58'h1;
  assign T32 = T23[3'h6:3'h6];
  assign T33 = T25[6'h3f:3'h6];
  assign io_replay = T34;
  assign T34 = io_host_ipi_req_valid & T35;
  assign T35 = io_host_ipi_req_ready ^ 1'h1;
  assign io_fatc = T36;
  assign T36 = wen & T37;
  assign T37 = T10[5'h11:5'h11];
  assign io_evec = T38;
  assign T38 = T39;
  assign T39 = io_exception ? T487 : reg_epc;
  assign T40 = T45 ? T43 : T41;
  assign T41 = io_exception ? T42 : reg_epc;
  assign T42 = io_pc;
  assign T43 = T44;
  assign T44 = wdata[6'h2b:1'h0];
  assign T45 = wen & T46;
  assign T46 = T10[3'h6:3'h6];
  assign T487 = {T488, T47};
  assign T47 = reg_evec;
  assign T48 = T51 ? T49 : reg_evec;
  assign T49 = T50;
  assign T50 = wdata[6'h2a:1'h0];
  assign T51 = wen & T52;
  assign T52 = T10[4'hc:4'hc];
  assign T488 = T47[6'h2a:6'h2a];
  assign io_ptbr = reg_ptbr;
  assign T53 = T57 ? T54 : reg_ptbr;
  assign T54 = T55;
  assign T55 = {T56, 13'h0};
  assign T56 = wdata[5'h1f:4'hd];
  assign T57 = wen & T58;
  assign T58 = T10[4'h8:4'h8];
  assign io_status_s = reg_status_s;
  assign T59 = reset ? 1'h1 : T60;
  assign T60 = T68 ? T67 : T61;
  assign T61 = io_sret ? reg_status_ps : T62;
  assign T62 = io_exception ? 1'h1 : reg_status_s;
  assign T63 = reset ? 1'h0 : T64;
  assign T64 = T68 ? T66 : T65;
  assign T65 = io_exception ? reg_status_s : reg_status_ps;
  assign T66 = wdata[1'h1:1'h1];
  assign T67 = wdata[1'h0:1'h0];
  assign T68 = wen & T69;
  assign T69 = T10[4'he:4'he];
  assign io_status_ps = reg_status_ps;
  assign io_status_ei = reg_status_ei;
  assign T70 = reset ? 1'h0 : T71;
  assign T71 = T68 ? T78 : T72;
  assign T72 = io_sret ? reg_status_pei : T73;
  assign T73 = io_exception ? 1'h0 : reg_status_ei;
  assign T74 = reset ? 1'h0 : T75;
  assign T75 = T68 ? T77 : T76;
  assign T76 = io_exception ? reg_status_ei : reg_status_pei;
  assign T77 = wdata[2'h3:2'h3];
  assign T78 = wdata[2'h2:2'h2];
  assign io_status_pei = reg_status_pei;
  assign io_status_ef = reg_status_ef;
  assign T79 = reset ? 1'h0 : T80;
  assign T80 = T68 ? T81 : reg_status_ef;
  assign T81 = wdata[3'h4:3'h4];
  assign io_status_u64 = reg_status_u64;
  assign T82 = reset ? 1'h1 : T83;
  assign T83 = T68 ? 1'h1 : T84;
  assign T84 = T68 ? T85 : reg_status_u64;
  assign T85 = wdata[3'h5:3'h5];
  assign io_status_s64 = reg_status_s64;
  assign T86 = reset ? 1'h1 : T87;
  assign T87 = T68 ? 1'h1 : T88;
  assign T88 = T68 ? T89 : reg_status_s64;
  assign T89 = wdata[3'h6:3'h6];
  assign io_status_vm = reg_status_vm;
  assign T90 = reset ? 1'h0 : T91;
  assign T91 = T68 ? T92 : reg_status_vm;
  assign T92 = wdata[3'h7:3'h7];
  assign io_status_er = reg_status_er;
  assign T93 = reset ? 1'h0 : T94;
  assign T94 = T68 ? 1'h0 : T95;
  assign T95 = T68 ? T96 : reg_status_er;
  assign T96 = wdata[4'h8:4'h8];
  assign io_status_zero = reg_status_zero;
  assign T97 = reset ? 7'h0 : T98;
  assign T98 = T68 ? 7'h0 : T99;
  assign T99 = T68 ? T100 : reg_status_zero;
  assign T100 = wdata[4'hf:4'h9];
  assign io_status_im = reg_status_im;
  assign T101 = reset ? 8'h0 : T102;
  assign T102 = T68 ? T103 : reg_status_im;
  assign T103 = wdata[5'h17:5'h10];
  assign io_status_ip = T104;
  assign T104 = {T105, 4'h0};
  assign T105 = {T112, T106};
  assign T106 = {r_irq_ipi, 1'h0};
  assign T489 = reset ? 1'h1 : T107;
  assign T107 = io_host_ipi_rep_valid ? 1'h1 : T108;
  assign T108 = T110 ? T109 : r_irq_ipi;
  assign T109 = wdata[1'h0:1'h0];
  assign T110 = wen & T111;
  assign T111 = T10[5'h13:5'h13];
  assign T112 = {r_irq_timer, T113};
  assign T113 = reg_fromhost != 64'h0;
  assign T490 = reset ? 64'h0 : T114;
  assign T114 = T115 ? wdata : reg_fromhost;
  assign T115 = T119 & T116;
  assign T116 = T118 | T117;
  assign T117 = host_pcr_req_fire ^ 1'h1;
  assign T118 = reg_fromhost == 64'h0;
  assign T119 = wen & T120;
  assign T120 = T10[5'h16:5'h16];
  assign T491 = reset ? 1'h0 : T121;
  assign T121 = T128 ? 1'h0 : T122;
  assign T122 = T123 ? 1'h1 : r_irq_timer;
  assign T123 = T127 == reg_compare;
  assign T124 = T128 ? T125 : reg_compare;
  assign T125 = T126;
  assign T126 = wdata[5'h1f:1'h0];
  assign T127 = T19[5'h1f:1'h0];
  assign T128 = wen & T129;
  assign T129 = T10[4'hb:4'hb];
  assign io_rw_rdata = T130;
  assign T130 = T144 | T131;
  assign T131 = T143 ? T132 : 64'h0;
  assign T132 = {R138, R133};
  assign T492 = reset ? 6'h0 : T134;
  assign T134 = T137 ? T135 : R133;
  assign T135 = T136[3'h5:1'h0];
  assign T136 = T493 + 7'h1;
  assign T493 = {1'h0, R133};
  assign T137 = io_uarch_counters_15 != 1'h0;
  assign T494 = reset ? 58'h0 : T139;
  assign T139 = T141 ? T140 : R138;
  assign T140 = R138 + 58'h1;
  assign T141 = T137 & T142;
  assign T142 = T136[3'h6:3'h6];
  assign T143 = T10[6'h2a:6'h2a];
  assign T144 = T158 | T145;
  assign T145 = T157 ? T146 : 64'h0;
  assign T146 = {R152, R147};
  assign T495 = reset ? 6'h0 : T148;
  assign T148 = T151 ? T149 : R147;
  assign T149 = T150[3'h5:1'h0];
  assign T150 = T496 + 7'h1;
  assign T496 = {1'h0, R147};
  assign T151 = io_uarch_counters_14 != 1'h0;
  assign T497 = reset ? 58'h0 : T153;
  assign T153 = T155 ? T154 : R152;
  assign T154 = R152 + 58'h1;
  assign T155 = T151 & T156;
  assign T156 = T150[3'h6:3'h6];
  assign T157 = T10[6'h29:6'h29];
  assign T158 = T172 | T159;
  assign T159 = T171 ? T160 : 64'h0;
  assign T160 = {R166, R161};
  assign T498 = reset ? 6'h0 : T162;
  assign T162 = T165 ? T163 : R161;
  assign T163 = T164[3'h5:1'h0];
  assign T164 = T499 + 7'h1;
  assign T499 = {1'h0, R161};
  assign T165 = io_uarch_counters_13 != 1'h0;
  assign T500 = reset ? 58'h0 : T167;
  assign T167 = T169 ? T168 : R166;
  assign T168 = R166 + 58'h1;
  assign T169 = T165 & T170;
  assign T170 = T164[3'h6:3'h6];
  assign T171 = T10[6'h28:6'h28];
  assign T172 = T186 | T173;
  assign T173 = T185 ? T174 : 64'h0;
  assign T174 = {R180, R175};
  assign T501 = reset ? 6'h0 : T176;
  assign T176 = T179 ? T177 : R175;
  assign T177 = T178[3'h5:1'h0];
  assign T178 = T502 + 7'h1;
  assign T502 = {1'h0, R175};
  assign T179 = io_uarch_counters_12 != 1'h0;
  assign T503 = reset ? 58'h0 : T181;
  assign T181 = T183 ? T182 : R180;
  assign T182 = R180 + 58'h1;
  assign T183 = T179 & T184;
  assign T184 = T178[3'h6:3'h6];
  assign T185 = T10[6'h27:6'h27];
  assign T186 = T200 | T187;
  assign T187 = T199 ? T188 : 64'h0;
  assign T188 = {R194, R189};
  assign T504 = reset ? 6'h0 : T190;
  assign T190 = T193 ? T191 : R189;
  assign T191 = T192[3'h5:1'h0];
  assign T192 = T505 + 7'h1;
  assign T505 = {1'h0, R189};
  assign T193 = io_uarch_counters_11 != 1'h0;
  assign T506 = reset ? 58'h0 : T195;
  assign T195 = T197 ? T196 : R194;
  assign T196 = R194 + 58'h1;
  assign T197 = T193 & T198;
  assign T198 = T192[3'h6:3'h6];
  assign T199 = T10[6'h26:6'h26];
  assign T200 = T214 | T201;
  assign T201 = T213 ? T202 : 64'h0;
  assign T202 = {R208, R203};
  assign T507 = reset ? 6'h0 : T204;
  assign T204 = T207 ? T205 : R203;
  assign T205 = T206[3'h5:1'h0];
  assign T206 = T508 + 7'h1;
  assign T508 = {1'h0, R203};
  assign T207 = io_uarch_counters_10 != 1'h0;
  assign T509 = reset ? 58'h0 : T209;
  assign T209 = T211 ? T210 : R208;
  assign T210 = R208 + 58'h1;
  assign T211 = T207 & T212;
  assign T212 = T206[3'h6:3'h6];
  assign T213 = T10[6'h25:6'h25];
  assign T214 = T228 | T215;
  assign T215 = T227 ? T216 : 64'h0;
  assign T216 = {R222, R217};
  assign T510 = reset ? 6'h0 : T218;
  assign T218 = T221 ? T219 : R217;
  assign T219 = T220[3'h5:1'h0];
  assign T220 = T511 + 7'h1;
  assign T511 = {1'h0, R217};
  assign T221 = io_uarch_counters_9 != 1'h0;
  assign T512 = reset ? 58'h0 : T223;
  assign T223 = T225 ? T224 : R222;
  assign T224 = R222 + 58'h1;
  assign T225 = T221 & T226;
  assign T226 = T220[3'h6:3'h6];
  assign T227 = T10[6'h24:6'h24];
  assign T228 = T242 | T229;
  assign T229 = T241 ? T230 : 64'h0;
  assign T230 = {R236, R231};
  assign T513 = reset ? 6'h0 : T232;
  assign T232 = T235 ? T233 : R231;
  assign T233 = T234[3'h5:1'h0];
  assign T234 = T514 + 7'h1;
  assign T514 = {1'h0, R231};
  assign T235 = io_uarch_counters_8 != 1'h0;
  assign T515 = reset ? 58'h0 : T237;
  assign T237 = T239 ? T238 : R236;
  assign T238 = R236 + 58'h1;
  assign T239 = T235 & T240;
  assign T240 = T234[3'h6:3'h6];
  assign T241 = T10[6'h23:6'h23];
  assign T242 = T256 | T243;
  assign T243 = T255 ? T244 : 64'h0;
  assign T244 = {R250, R245};
  assign T516 = reset ? 6'h0 : T246;
  assign T246 = T249 ? T247 : R245;
  assign T247 = T248[3'h5:1'h0];
  assign T248 = T517 + 7'h1;
  assign T517 = {1'h0, R245};
  assign T249 = io_uarch_counters_7 != 1'h0;
  assign T518 = reset ? 58'h0 : T251;
  assign T251 = T253 ? T252 : R250;
  assign T252 = R250 + 58'h1;
  assign T253 = T249 & T254;
  assign T254 = T248[3'h6:3'h6];
  assign T255 = T10[6'h22:6'h22];
  assign T256 = T270 | T257;
  assign T257 = T269 ? T258 : 64'h0;
  assign T258 = {R264, R259};
  assign T519 = reset ? 6'h0 : T260;
  assign T260 = T263 ? T261 : R259;
  assign T261 = T262[3'h5:1'h0];
  assign T262 = T520 + 7'h1;
  assign T520 = {1'h0, R259};
  assign T263 = io_uarch_counters_6 != 1'h0;
  assign T521 = reset ? 58'h0 : T265;
  assign T265 = T267 ? T266 : R264;
  assign T266 = R264 + 58'h1;
  assign T267 = T263 & T268;
  assign T268 = T262[3'h6:3'h6];
  assign T269 = T10[6'h21:6'h21];
  assign T270 = T284 | T271;
  assign T271 = T283 ? T272 : 64'h0;
  assign T272 = {R278, R273};
  assign T522 = reset ? 6'h0 : T274;
  assign T274 = T277 ? T275 : R273;
  assign T275 = T276[3'h5:1'h0];
  assign T276 = T523 + 7'h1;
  assign T523 = {1'h0, R273};
  assign T277 = io_uarch_counters_5 != 1'h0;
  assign T524 = reset ? 58'h0 : T279;
  assign T279 = T281 ? T280 : R278;
  assign T280 = R278 + 58'h1;
  assign T281 = T277 & T282;
  assign T282 = T276[3'h6:3'h6];
  assign T283 = T10[6'h20:6'h20];
  assign T284 = T298 | T285;
  assign T285 = T297 ? T286 : 64'h0;
  assign T286 = {R292, R287};
  assign T525 = reset ? 6'h0 : T288;
  assign T288 = T291 ? T289 : R287;
  assign T289 = T290[3'h5:1'h0];
  assign T290 = T526 + 7'h1;
  assign T526 = {1'h0, R287};
  assign T291 = io_uarch_counters_4 != 1'h0;
  assign T527 = reset ? 58'h0 : T293;
  assign T293 = T295 ? T294 : R292;
  assign T294 = R292 + 58'h1;
  assign T295 = T291 & T296;
  assign T296 = T290[3'h6:3'h6];
  assign T297 = T10[5'h1f:5'h1f];
  assign T298 = T312 | T299;
  assign T299 = T311 ? T300 : 64'h0;
  assign T300 = {R306, R301};
  assign T528 = reset ? 6'h0 : T302;
  assign T302 = T305 ? T303 : R301;
  assign T303 = T304[3'h5:1'h0];
  assign T304 = T529 + 7'h1;
  assign T529 = {1'h0, R301};
  assign T305 = io_uarch_counters_3 != 1'h0;
  assign T530 = reset ? 58'h0 : T307;
  assign T307 = T309 ? T308 : R306;
  assign T308 = R306 + 58'h1;
  assign T309 = T305 & T310;
  assign T310 = T304[3'h6:3'h6];
  assign T311 = T10[5'h1e:5'h1e];
  assign T312 = T326 | T313;
  assign T313 = T325 ? T314 : 64'h0;
  assign T314 = {R320, R315};
  assign T531 = reset ? 6'h0 : T316;
  assign T316 = T319 ? T317 : R315;
  assign T317 = T318[3'h5:1'h0];
  assign T318 = T532 + 7'h1;
  assign T532 = {1'h0, R315};
  assign T319 = io_uarch_counters_2 != 1'h0;
  assign T533 = reset ? 58'h0 : T321;
  assign T321 = T323 ? T322 : R320;
  assign T322 = R320 + 58'h1;
  assign T323 = T319 & T324;
  assign T324 = T318[3'h6:3'h6];
  assign T325 = T10[5'h1d:5'h1d];
  assign T326 = T340 | T327;
  assign T327 = T339 ? T328 : 64'h0;
  assign T328 = {R334, R329};
  assign T534 = reset ? 6'h0 : T330;
  assign T330 = T333 ? T331 : R329;
  assign T331 = T332[3'h5:1'h0];
  assign T332 = T535 + 7'h1;
  assign T535 = {1'h0, R329};
  assign T333 = io_uarch_counters_1 != 1'h0;
  assign T536 = reset ? 58'h0 : T335;
  assign T335 = T337 ? T336 : R334;
  assign T336 = R334 + 58'h1;
  assign T337 = T333 & T338;
  assign T338 = T332[3'h6:3'h6];
  assign T339 = T10[5'h1c:5'h1c];
  assign T340 = T354 | T341;
  assign T341 = T353 ? T342 : 64'h0;
  assign T342 = {R348, R343};
  assign T537 = reset ? 6'h0 : T344;
  assign T344 = T347 ? T345 : R343;
  assign T345 = T346[3'h5:1'h0];
  assign T346 = T538 + 7'h1;
  assign T538 = {1'h0, R343};
  assign T347 = io_uarch_counters_0 != 1'h0;
  assign T539 = reset ? 58'h0 : T349;
  assign T349 = T351 ? T350 : R348;
  assign T350 = R348 + 58'h1;
  assign T351 = T347 & T352;
  assign T352 = T346[3'h6:3'h6];
  assign T353 = T10[5'h1b:5'h1b];
  assign T354 = T356 | T355;
  assign T355 = T120 ? reg_fromhost : 64'h0;
  assign T356 = T368 | T357;
  assign T357 = T367 ? reg_tohost : 64'h0;
  assign T540 = reset ? 64'h0 : T358;
  assign T358 = T363 ? wdata : T359;
  assign T359 = T360 ? 64'h0 : reg_tohost;
  assign T360 = T361 & T367;
  assign T361 = host_pcr_req_fire & T362;
  assign T362 = host_pcr_bits_rw ^ 1'h1;
  assign T363 = T366 & T364;
  assign T364 = T365 | host_pcr_req_fire;
  assign T365 = reg_tohost == 64'h0;
  assign T366 = wen & T367;
  assign T367 = T10[5'h15:5'h15];
  assign T368 = T374 | T541;
  assign T541 = {63'h0, T369};
  assign T369 = T373 ? reg_stats : 1'h0;
  assign T542 = reset ? 1'h0 : T370;
  assign T370 = T372 ? T371 : reg_stats;
  assign T371 = wdata[1'h0:1'h0];
  assign T372 = wen & T373;
  assign T373 = T10[2'h3:2'h3];
  assign T374 = T376 | T543;
  assign T543 = {62'h0, T375};
  assign T375 = T111 ? 2'h2 : 2'h0;
  assign T376 = T379 | T544;
  assign T544 = {62'h0, T377};
  assign T377 = T378 ? 2'h2 : 2'h0;
  assign T378 = T10[5'h12:5'h12];
  assign T379 = T381 | T545;
  assign T545 = {62'h0, T380};
  assign T380 = T37 ? 2'h2 : 2'h0;
  assign T381 = T384 | T546;
  assign T546 = {62'h0, T382};
  assign T382 = T383 ? 2'h2 : 2'h0;
  assign T383 = T10[5'h10:5'h10];
  assign T384 = T387 | T547;
  assign T547 = {63'h0, T385};
  assign T385 = T386 ? io_host_id : 1'h0;
  assign T386 = T10[4'hf:4'hf];
  assign T387 = T401 | T548;
  assign T548 = {32'h0, T388};
  assign T388 = T69 ? T389 : 32'h0;
  assign T389 = T390;
  assign T390 = {T396, T391};
  assign T391 = {T394, T392};
  assign T392 = {io_status_ei, T393};
  assign T393 = {io_status_ps, io_status_s};
  assign T394 = {io_status_u64, T395};
  assign T395 = {io_status_ef, io_status_pei};
  assign T396 = {T399, T397};
  assign T397 = {io_status_er, T398};
  assign T398 = {io_status_vm, io_status_s64};
  assign T399 = {io_status_ip, T400};
  assign T400 = {io_status_im, io_status_zero};
  assign T401 = T405 | T402;
  assign T402 = T404 ? reg_cause : 64'h0;
  assign T403 = io_exception ? io_cause : reg_cause;
  assign T404 = T10[4'hd:4'hd];
  assign T405 = T407 | T549;
  assign T549 = {21'h0, T406};
  assign T406 = T52 ? reg_evec : 43'h0;
  assign T407 = T409 | T550;
  assign T550 = {32'h0, T408};
  assign T408 = T129 ? reg_compare : 32'h0;
  assign T409 = T411 | T410;
  assign T410 = T27 ? T19 : 64'h0;
  assign T411 = T412 | 64'h0;
  assign T412 = T415 | T551;
  assign T551 = {32'h0, T413};
  assign T413 = T58 ? read_ptbr : 32'h0;
  assign read_ptbr = T414 << 4'hd;
  assign T414 = reg_ptbr[5'h1f:4'hd];
  assign T415 = T428 | T552;
  assign T552 = {21'h0, T416};
  assign T416 = T427 ? reg_badvaddr : 43'h0;
  assign T553 = T417[6'h2a:1'h0];
  assign T417 = io_badvaddr_wen ? T418 : T554;
  assign T554 = {1'h0, reg_badvaddr};
  assign T418 = T419;
  assign T419 = {T421, T420};
  assign T420 = io_rw_wdata[6'h2a:1'h0];
  assign T421 = T425 ? T424 : T422;
  assign T422 = T423 != 21'h0;
  assign T423 = io_rw_wdata[6'h3f:6'h2b];
  assign T424 = T423 == 21'h1fffff;
  assign T425 = $signed(T426) < $signed(1'h0);
  assign T426 = T420;
  assign T427 = T10[3'h7:3'h7];
  assign T428 = T430 | T555;
  assign T555 = {20'h0, T429};
  assign T429 = T46 ? reg_epc : 44'h0;
  assign T430 = T435 | T431;
  assign T431 = T434 ? reg_sup1 : 64'h0;
  assign T432 = T433 ? wdata : reg_sup1;
  assign T433 = wen & T434;
  assign T434 = T10[3'h5:3'h5];
  assign T435 = T440 | T436;
  assign T436 = T439 ? reg_sup0 : 64'h0;
  assign T437 = T438 ? wdata : reg_sup0;
  assign T438 = wen & T439;
  assign T439 = T10[3'h4:3'h4];
  assign T440 = T454 | T441;
  assign T441 = T453 ? T442 : 64'h0;
  assign T442 = {R448, R443};
  assign T556 = reset ? 6'h0 : T444;
  assign T444 = T447 ? T445 : R443;
  assign T445 = T446[3'h5:1'h0];
  assign T446 = T557 + 7'h1;
  assign T557 = {1'h0, R443};
  assign T447 = io_retire != 1'h0;
  assign T558 = reset ? 58'h0 : T449;
  assign T449 = T451 ? T450 : R448;
  assign T450 = R448 + 58'h1;
  assign T451 = T447 & T452;
  assign T452 = T446[3'h6:3'h6];
  assign T453 = T10[5'h1a:5'h1a];
  assign T454 = T457 | T455;
  assign T455 = T456 ? T19 : 64'h0;
  assign T456 = T10[5'h19:5'h19];
  assign T457 = T559 | T458;
  assign T458 = T459 ? T19 : 64'h0;
  assign T459 = T10[5'h18:5'h18];
  assign T559 = {56'h0, T460};
  assign T460 = T562 | T461;
  assign T461 = T18 ? T462 : 8'h0;
  assign T462 = {reg_frm, reg_fflags};
  assign T560 = T463[3'h4:1'h0];
  assign T463 = T17 ? wdata : T464;
  assign T464 = T467 ? wdata : T561;
  assign T561 = {59'h0, T465};
  assign T465 = io_fcsr_flags_valid ? T466 : reg_fflags;
  assign T466 = reg_fflags | io_fcsr_flags_bits;
  assign T467 = wen & T468;
  assign T468 = T10[1'h0:1'h0];
  assign T562 = {3'h0, T469};
  assign T469 = T471 | T563;
  assign T563 = {2'h0, T470};
  assign T470 = T9 ? reg_frm : 3'h0;
  assign T471 = T468 ? reg_fflags : 5'h0;
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T564;
  assign T564 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T472;
  assign T472 = cpu_req_valid & T378;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T473 = T475 ? 1'h0 : T474;
  assign T474 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T475 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T476;
  assign T476 = T478 & T477;
  assign T477 = host_pcr_rep_valid ^ 1'h1;
  assign T478 = host_pcr_req_valid ^ 1'h1;

  always @(posedge clk) begin
    reg_frm <= T479;
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T4) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T4) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(T4) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T4) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    if(reset) begin
      R20 <= 6'h0;
    end else if(T26) begin
      R20 <= T24;
    end else begin
      R20 <= T22;
    end
    if(reset) begin
      R28 <= 58'h0;
    end else if(T26) begin
      R28 <= T33;
    end else if(T32) begin
      R28 <= T31;
    end
    if(T45) begin
      reg_epc <= T43;
    end else if(io_exception) begin
      reg_epc <= T42;
    end
    if(T51) begin
      reg_evec <= T49;
    end
    if(T57) begin
      reg_ptbr <= T54;
    end
    if(reset) begin
      reg_status_s <= 1'h1;
    end else if(T68) begin
      reg_status_s <= T67;
    end else if(io_sret) begin
      reg_status_s <= reg_status_ps;
    end else if(io_exception) begin
      reg_status_s <= 1'h1;
    end
    if(reset) begin
      reg_status_ps <= 1'h0;
    end else if(T68) begin
      reg_status_ps <= T66;
    end else if(io_exception) begin
      reg_status_ps <= reg_status_s;
    end
    if(reset) begin
      reg_status_ei <= 1'h0;
    end else if(T68) begin
      reg_status_ei <= T78;
    end else if(io_sret) begin
      reg_status_ei <= reg_status_pei;
    end else if(io_exception) begin
      reg_status_ei <= 1'h0;
    end
    if(reset) begin
      reg_status_pei <= 1'h0;
    end else if(T68) begin
      reg_status_pei <= T77;
    end else if(io_exception) begin
      reg_status_pei <= reg_status_ei;
    end
    if(reset) begin
      reg_status_ef <= 1'h0;
    end else if(T68) begin
      reg_status_ef <= T81;
    end
    if(reset) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= T85;
    end
    if(reset) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= T89;
    end
    if(reset) begin
      reg_status_vm <= 1'h0;
    end else if(T68) begin
      reg_status_vm <= T92;
    end
    if(reset) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= T96;
    end
    if(reset) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= T100;
    end
    if(reset) begin
      reg_status_im <= 8'h0;
    end else if(T68) begin
      reg_status_im <= T103;
    end
    if(reset) begin
      r_irq_ipi <= 1'h1;
    end else if(io_host_ipi_rep_valid) begin
      r_irq_ipi <= 1'h1;
    end else if(T110) begin
      r_irq_ipi <= T109;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T115) begin
      reg_fromhost <= wdata;
    end
    if(reset) begin
      r_irq_timer <= 1'h0;
    end else if(T128) begin
      r_irq_timer <= 1'h0;
    end else if(T123) begin
      r_irq_timer <= 1'h1;
    end
    if(T128) begin
      reg_compare <= T125;
    end
    if(reset) begin
      R133 <= 6'h0;
    end else if(T137) begin
      R133 <= T135;
    end
    if(reset) begin
      R138 <= 58'h0;
    end else if(T141) begin
      R138 <= T140;
    end
    if(reset) begin
      R147 <= 6'h0;
    end else if(T151) begin
      R147 <= T149;
    end
    if(reset) begin
      R152 <= 58'h0;
    end else if(T155) begin
      R152 <= T154;
    end
    if(reset) begin
      R161 <= 6'h0;
    end else if(T165) begin
      R161 <= T163;
    end
    if(reset) begin
      R166 <= 58'h0;
    end else if(T169) begin
      R166 <= T168;
    end
    if(reset) begin
      R175 <= 6'h0;
    end else if(T179) begin
      R175 <= T177;
    end
    if(reset) begin
      R180 <= 58'h0;
    end else if(T183) begin
      R180 <= T182;
    end
    if(reset) begin
      R189 <= 6'h0;
    end else if(T193) begin
      R189 <= T191;
    end
    if(reset) begin
      R194 <= 58'h0;
    end else if(T197) begin
      R194 <= T196;
    end
    if(reset) begin
      R203 <= 6'h0;
    end else if(T207) begin
      R203 <= T205;
    end
    if(reset) begin
      R208 <= 58'h0;
    end else if(T211) begin
      R208 <= T210;
    end
    if(reset) begin
      R217 <= 6'h0;
    end else if(T221) begin
      R217 <= T219;
    end
    if(reset) begin
      R222 <= 58'h0;
    end else if(T225) begin
      R222 <= T224;
    end
    if(reset) begin
      R231 <= 6'h0;
    end else if(T235) begin
      R231 <= T233;
    end
    if(reset) begin
      R236 <= 58'h0;
    end else if(T239) begin
      R236 <= T238;
    end
    if(reset) begin
      R245 <= 6'h0;
    end else if(T249) begin
      R245 <= T247;
    end
    if(reset) begin
      R250 <= 58'h0;
    end else if(T253) begin
      R250 <= T252;
    end
    if(reset) begin
      R259 <= 6'h0;
    end else if(T263) begin
      R259 <= T261;
    end
    if(reset) begin
      R264 <= 58'h0;
    end else if(T267) begin
      R264 <= T266;
    end
    if(reset) begin
      R273 <= 6'h0;
    end else if(T277) begin
      R273 <= T275;
    end
    if(reset) begin
      R278 <= 58'h0;
    end else if(T281) begin
      R278 <= T280;
    end
    if(reset) begin
      R287 <= 6'h0;
    end else if(T291) begin
      R287 <= T289;
    end
    if(reset) begin
      R292 <= 58'h0;
    end else if(T295) begin
      R292 <= T294;
    end
    if(reset) begin
      R301 <= 6'h0;
    end else if(T305) begin
      R301 <= T303;
    end
    if(reset) begin
      R306 <= 58'h0;
    end else if(T309) begin
      R306 <= T308;
    end
    if(reset) begin
      R315 <= 6'h0;
    end else if(T319) begin
      R315 <= T317;
    end
    if(reset) begin
      R320 <= 58'h0;
    end else if(T323) begin
      R320 <= T322;
    end
    if(reset) begin
      R329 <= 6'h0;
    end else if(T333) begin
      R329 <= T331;
    end
    if(reset) begin
      R334 <= 58'h0;
    end else if(T337) begin
      R334 <= T336;
    end
    if(reset) begin
      R343 <= 6'h0;
    end else if(T347) begin
      R343 <= T345;
    end
    if(reset) begin
      R348 <= 58'h0;
    end else if(T351) begin
      R348 <= T350;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T363) begin
      reg_tohost <= wdata;
    end else if(T360) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T372) begin
      reg_stats <= T371;
    end
    if(io_exception) begin
      reg_cause <= io_cause;
    end
    reg_badvaddr <= T553;
    if(T433) begin
      reg_sup1 <= wdata;
    end
    if(T438) begin
      reg_sup0 <= wdata;
    end
    if(reset) begin
      R443 <= 6'h0;
    end else if(T447) begin
      R443 <= T445;
    end
    if(reset) begin
      R448 <= 58'h0;
    end else if(T451) begin
      R448 <= T450;
    end
    reg_fflags <= T560;
    if(T475) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module Datapath(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [2:0] io_ctrl_sel_pc,
    input  io_ctrl_killd,
    input  io_ctrl_killm,
    input  io_ctrl_ren_1,
    input  io_ctrl_ren_0,
    input  io_ctrl_ex_ctrl_legal,
    input  io_ctrl_ex_ctrl_fp,
    input  io_ctrl_ex_ctrl_rocc,
    input  io_ctrl_ex_ctrl_branch,
    input  io_ctrl_ex_ctrl_jal,
    input  io_ctrl_ex_ctrl_jalr,
    input  io_ctrl_ex_ctrl_rxs2,
    input  io_ctrl_ex_ctrl_rxs1,
    input [1:0] io_ctrl_ex_ctrl_sel_alu2,
    input [1:0] io_ctrl_ex_ctrl_sel_alu1,
    input [2:0] io_ctrl_ex_ctrl_sel_imm,
    input  io_ctrl_ex_ctrl_alu_dw,
    input [3:0] io_ctrl_ex_ctrl_alu_fn,
    input  io_ctrl_ex_ctrl_mem,
    input [4:0] io_ctrl_ex_ctrl_mem_cmd,
    input [3:0] io_ctrl_ex_ctrl_mem_type,
    input  io_ctrl_ex_ctrl_rfs1,
    input  io_ctrl_ex_ctrl_rfs2,
    input  io_ctrl_ex_ctrl_rfs3,
    input  io_ctrl_ex_ctrl_wfd,
    input  io_ctrl_ex_ctrl_div,
    input  io_ctrl_ex_ctrl_wxd,
    input [1:0] io_ctrl_ex_ctrl_csr,
    input  io_ctrl_ex_ctrl_fence_i,
    input  io_ctrl_ex_ctrl_sret,
    input  io_ctrl_ex_ctrl_scall,
    input  io_ctrl_ex_ctrl_fence,
    input  io_ctrl_ex_ctrl_amo,
    input  io_ctrl_mem_ctrl_legal,
    input  io_ctrl_mem_ctrl_fp,
    input  io_ctrl_mem_ctrl_rocc,
    input  io_ctrl_mem_ctrl_branch,
    input  io_ctrl_mem_ctrl_jal,
    input  io_ctrl_mem_ctrl_jalr,
    input  io_ctrl_mem_ctrl_rxs2,
    input  io_ctrl_mem_ctrl_rxs1,
    input [1:0] io_ctrl_mem_ctrl_sel_alu2,
    input [1:0] io_ctrl_mem_ctrl_sel_alu1,
    input [2:0] io_ctrl_mem_ctrl_sel_imm,
    input  io_ctrl_mem_ctrl_alu_dw,
    input [3:0] io_ctrl_mem_ctrl_alu_fn,
    input  io_ctrl_mem_ctrl_mem,
    input [4:0] io_ctrl_mem_ctrl_mem_cmd,
    input [3:0] io_ctrl_mem_ctrl_mem_type,
    input  io_ctrl_mem_ctrl_rfs1,
    input  io_ctrl_mem_ctrl_rfs2,
    input  io_ctrl_mem_ctrl_rfs3,
    input  io_ctrl_mem_ctrl_wfd,
    input  io_ctrl_mem_ctrl_div,
    input  io_ctrl_mem_ctrl_wxd,
    input [1:0] io_ctrl_mem_ctrl_csr,
    input  io_ctrl_mem_ctrl_fence_i,
    input  io_ctrl_mem_ctrl_sret,
    input  io_ctrl_mem_ctrl_scall,
    input  io_ctrl_mem_ctrl_fence,
    input  io_ctrl_mem_ctrl_amo,
    input [2:0] io_ctrl_csr,
    input  io_ctrl_sret,
    input  io_ctrl_ex_valid,
    input  io_ctrl_wb_wen,
    input  io_ctrl_bypass_1,
    input  io_ctrl_bypass_0,
    input [1:0] io_ctrl_bypass_src_1,
    input [1:0] io_ctrl_bypass_src_0,
    input  io_ctrl_ll_ready,
    input  io_ctrl_retire,
    input  io_ctrl_exception,
    input [63:0] io_ctrl_cause,
    input  io_ctrl_badvaddr_wen,
    output[31:0] io_ctrl_inst,
    output io_ctrl_mem_br_taken,
    output io_ctrl_mem_misprediction,
    output io_ctrl_div_mul_rdy,
    output io_ctrl_ll_wen,
    output[4:0] io_ctrl_ll_waddr,
    output[4:0] io_ctrl_ex_waddr,
    output io_ctrl_mem_rs1_ra,
    output[4:0] io_ctrl_mem_waddr,
    output[4:0] io_ctrl_wb_waddr,
    output[7:0] io_ctrl_status_ip,
    output[7:0] io_ctrl_status_im,
    output[6:0] io_ctrl_status_zero,
    output io_ctrl_status_er,
    output io_ctrl_status_vm,
    output io_ctrl_status_s64,
    output io_ctrl_status_u64,
    output io_ctrl_status_ef,
    output io_ctrl_status_pei,
    output io_ctrl_status_ei,
    output io_ctrl_status_ps,
    output io_ctrl_status_s,
    output io_ctrl_fp_sboard_clr,
    output[4:0] io_ctrl_fp_sboard_clra,
    output io_ctrl_csr_replay,
    input  io_dmem_req_ready,
    //output io_dmem_req_valid
    //output io_dmem_req_bits_kill
    //output[3:0] io_dmem_req_bits_typ
    //output io_dmem_req_bits_phys
    output[43:0] io_dmem_req_bits_addr,
    output[7:0] io_dmem_req_bits_tag,
    //output[4:0] io_dmem_req_bits_cmd
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [3:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    //output io_imem_req_valid
    output[43:0] io_imem_req_bits_pc,
    //output io_imem_resp_ready
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    //output io_imem_btb_update_valid
    //output io_imem_btb_update_bits_prediction_valid
    //output io_imem_btb_update_bits_prediction_bits_taken
    //output io_imem_btb_update_bits_prediction_bits_mask
    //output io_imem_btb_update_bits_prediction_bits_bridx
    //output[42:0] io_imem_btb_update_bits_prediction_bits_target
    //output[5:0] io_imem_btb_update_bits_prediction_bits_entry
    //output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history
    //output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    //output io_imem_btb_update_bits_taken
    //output io_imem_btb_update_bits_isJump
    //output io_imem_btb_update_bits_isReturn
    output[42:0] io_imem_btb_update_bits_br_pc,
    //output io_imem_bht_update_valid
    //output io_imem_bht_update_bits_prediction_valid
    //output io_imem_bht_update_bits_prediction_bits_taken
    //output io_imem_bht_update_bits_prediction_bits_mask
    //output io_imem_bht_update_bits_prediction_bits_bridx
    //output[42:0] io_imem_bht_update_bits_prediction_bits_target
    //output[5:0] io_imem_bht_update_bits_prediction_bits_entry
    //output[6:0] io_imem_bht_update_bits_prediction_bits_bht_history
    //output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_bht_update_bits_pc,
    //output io_imem_bht_update_bits_taken
    //output io_imem_bht_update_bits_mispredict
    //output io_imem_ras_update_valid
    //output io_imem_ras_update_bits_isCall
    //output io_imem_ras_update_bits_isReturn
    output[42:0] io_imem_ras_update_bits_returnAddr,
    //output io_imem_ras_update_bits_prediction_valid
    //output io_imem_ras_update_bits_prediction_bits_taken
    //output io_imem_ras_update_bits_prediction_bits_mask
    //output io_imem_ras_update_bits_prediction_bits_bridx
    //output[42:0] io_imem_ras_update_bits_prediction_bits_target
    //output[5:0] io_imem_ras_update_bits_prediction_bits_entry
    //output[6:0] io_imem_ras_update_bits_prediction_bits_bht_history
    //output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    //output io_imem_invalidate
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [3:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[3:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[135:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_manager_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_manager_xact_id,
    //output io_rocc_dmem_acquire_ready
    input  io_rocc_dmem_acquire_valid,
    input [1:0] io_rocc_dmem_acquire_bits_header_src,
    input [1:0] io_rocc_dmem_acquire_bits_header_dst,
    input [25:0] io_rocc_dmem_acquire_bits_payload_addr,
    input [1:0] io_rocc_dmem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_acquire_bits_payload_data,
    input  io_rocc_dmem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_dmem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_dmem_acquire_bits_payload_subblock,
    input  io_rocc_dmem_grant_ready,
    //output io_rocc_dmem_grant_valid
    //output[1:0] io_rocc_dmem_grant_bits_header_src
    //output[1:0] io_rocc_dmem_grant_bits_header_dst
    //output[135:0] io_rocc_dmem_grant_bits_payload_data
    //output[1:0] io_rocc_dmem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_dmem_grant_bits_payload_manager_xact_id
    //output io_rocc_dmem_grant_bits_payload_uncached
    //output[1:0] io_rocc_dmem_grant_bits_payload_g_type
    //output io_rocc_dmem_finish_ready
    input  io_rocc_dmem_finish_valid,
    input [1:0] io_rocc_dmem_finish_bits_header_src,
    input [1:0] io_rocc_dmem_finish_bits_header_dst,
    input [3:0] io_rocc_dmem_finish_bits_payload_manager_xact_id,
    input  io_rocc_dmem_probe_ready,
    //output io_rocc_dmem_probe_valid
    //output[1:0] io_rocc_dmem_probe_bits_header_src
    //output[1:0] io_rocc_dmem_probe_bits_header_dst
    //output[25:0] io_rocc_dmem_probe_bits_payload_addr
    //output[1:0] io_rocc_dmem_probe_bits_payload_p_type
    //output io_rocc_dmem_release_ready
    input  io_rocc_dmem_release_valid,
    input [1:0] io_rocc_dmem_release_bits_header_src,
    input [1:0] io_rocc_dmem_release_bits_header_dst,
    input [25:0] io_rocc_dmem_release_bits_payload_addr,
    input [1:0] io_rocc_dmem_release_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_release_bits_payload_data,
    input [2:0] io_rocc_dmem_release_bits_payload_r_type,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  reg  ex_reg_kill;
  wire T7;
  reg  mem_reg_kill;
  wire[31:0] T8;
  wire[63:0] T9;
  reg [63:0] R10;
  reg [63:0] R11;
  wire[63:0] ex_rs_1;
  wire[63:0] T12;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[63:0] id_rs_1;
  wire[63:0] T16;
  wire[63:0] T17;
  reg [63:0] T18 [30:0];
  wire[63:0] T19;
  wire T20;
  wire T21;
  wire[4:0] T22;
  wire T23;
  wire T24;
  wire[4:0] wb_waddr;
  wire wb_wen;
  wire[4:0] T25;
  wire[4:0] T26;
  wire[4:0] T27;
  wire[63:0] wb_wdata;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  reg [63:0] wb_reg_wdata;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] mem_int_wdata;
  reg [63:0] mem_reg_wdata;
  wire[63:0] T33;
  wire[63:0] T281;
  wire[44:0] mem_br_target;
  wire[44:0] T34;
  wire[44:0] T35;
  reg [43:0] mem_reg_pc;
  wire[43:0] T36;
  reg [43:0] ex_reg_pc;
  wire[43:0] T37;
  wire[44:0] T282;
  wire[21:0] T38;
  wire[21:0] T39;
  wire[21:0] T40;
  wire[21:0] T41;
  wire[11:0] T42;
  wire[4:0] T43;
  wire[3:0] T44;
  wire[6:0] T45;
  wire[5:0] T46;
  wire T47;
  wire T48;
  wire[9:0] T49;
  wire[8:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire T53;
  wire T54;
  wire[21:0] T283;
  wire[14:0] T55;
  wire[14:0] T56;
  wire[11:0] T57;
  wire[4:0] T58;
  wire[3:0] T59;
  wire[6:0] T60;
  wire[5:0] T61;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire[1:0] T65;
  wire T66;
  wire T67;
  wire[6:0] T284;
  wire T285;
  wire T68;
  wire[22:0] T286;
  wire T287;
  wire[18:0] T288;
  wire T289;
  wire T69;
  wire T70;
  wire[63:0] ll_wdata;
  wire T71;
  wire dmem_resp_xpu;
  wire T72;
  wire T73;
  wire dmem_resp_valid;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T78;
  wire[61:0] T79;
  wire T80;
  wire T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[63:0] T290;
  wire bypass_0;
  wire[63:0] bypass_1;
  wire T84;
  wire[1:0] T85;
  wire[63:0] T86;
  wire[63:0] bypass_2;
  wire[63:0] bypass_3;
  wire T87;
  wire T88;
  reg  ex_reg_rs_bypass_1;
  wire T89;
  wire[4:0] T90;
  wire[4:0] T91;
  wire[63:0] T92;
  reg [63:0] R93;
  reg [63:0] R94;
  wire[63:0] ex_rs_0;
  wire[63:0] T95;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire[63:0] id_rs_0;
  wire[63:0] T99;
  wire[63:0] T100;
  wire[4:0] T101;
  wire[4:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T107;
  wire[61:0] T108;
  wire T109;
  wire T110;
  wire[63:0] T111;
  wire[63:0] T112;
  wire[63:0] T291;
  wire T113;
  wire[1:0] T114;
  wire[63:0] T115;
  wire T116;
  wire T117;
  reg  ex_reg_rs_bypass_0;
  wire T118;
  wire[4:0] T119;
  wire[4:0] T120;
  wire T121;
  wire[63:0] T122;
  wire[4:0] T123;
  wire[4:0] T124;
  wire[43:0] T125;
  reg [43:0] wb_reg_pc;
  wire[43:0] T126;
  wire T127;
  wire[32:0] T128;
  wire[32:0] T129;
  wire T130;
  wire[1135:0] T131;
  wire[63:0] T132;
  wire[63:0] T133;
  wire[63:0] T134;
  wire[63:0] T135;
  wire T136;
  wire[63:0] T137;
  wire T138;
  wire[1:0] T292;
  wire[11:0] T139;
  wire T140;
  wire T141;
  wire dmem_resp_replay;
  wire T142;
  reg  R143;
  wire T144;
  wire T145;
  wire[63:0] ex_op1;
  wire[63:0] T293;
  wire[43:0] T146;
  wire[43:0] T147;
  wire T148;
  wire[19:0] T294;
  wire T295;
  wire[63:0] T149;
  wire T150;
  wire[63:0] T151;
  wire[63:0] ex_op2;
  wire[63:0] T296;
  wire[31:0] T152;
  wire[31:0] T297;
  wire[3:0] T153;
  wire T154;
  wire[27:0] T298;
  wire T299;
  wire[31:0] ex_imm;
  wire[31:0] T155;
  wire[11:0] T156;
  wire[4:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire[3:0] T167;
  wire[3:0] T168;
  wire[3:0] T169;
  wire[3:0] T170;
  wire[3:0] T171;
  wire T172;
  wire[3:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire[6:0] T178;
  wire[5:0] T179;
  wire[5:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[19:0] T198;
  wire[18:0] T199;
  wire[7:0] T200;
  wire[7:0] T201;
  wire[7:0] T202;
  wire[7:0] T300;
  wire T203;
  wire T204;
  wire T205;
  wire[10:0] T206;
  wire[10:0] T301;
  wire[10:0] T207;
  wire[10:0] T208;
  wire T209;
  wire T210;
  wire[31:0] T302;
  wire T303;
  wire[63:0] T211;
  wire T212;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T213;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire[6:0] T219;
  wire[4:0] T220;
  wire T221;
  wire T222;
  wire T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[6:0] T226;
  wire[4:0] T304;
  wire[6:0] dmem_resp_waddr;
  wire[7:0] T227;
  wire[2:0] T305;
  wire T228;
  wire dmem_resp_fpu;
  wire T229;
  wire[42:0] T306;
  wire[42:0] T307;
  wire[42:0] T308;
  wire[42:0] T309;
  wire[42:0] T310;
  wire[43:0] T311;
  wire[44:0] T230;
  wire[44:0] T231;
  wire[44:0] T312;
  wire[43:0] T232;
  wire T233;
  wire[44:0] mem_npc;
  wire[44:0] T313;
  wire[43:0] T234;
  wire[42:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire[1:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[21:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire[63:0] T250;
  wire[7:0] T314;
  wire[5:0] T251;
  wire[43:0] T252;
  wire[43:0] T253;
  wire[42:0] T254;
  wire T255;
  wire T256;
  wire T257;
  wire[1:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire[21:0] T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[4:0] T315;
  wire T268;
  wire[4:0] T269;
  wire[4:0] T270;
  wire T271;
  wire[4:0] T272;
  wire[4:0] T273;
  wire[4:0] T316;
  wire[6:0] T274;
  wire[6:0] T317;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[44:0] T318;
  wire T280;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;
  wire pcr_io_host_pcr_req_ready;
  wire pcr_io_host_pcr_rep_valid;
  wire[63:0] pcr_io_host_pcr_rep_bits;
  wire pcr_io_host_ipi_req_valid;
  wire pcr_io_host_ipi_req_bits;
  wire pcr_io_host_ipi_rep_ready;
  wire pcr_io_host_debug_stats_pcr;
  wire[63:0] pcr_io_rw_rdata;
  wire[7:0] pcr_io_status_ip;
  wire[7:0] pcr_io_status_im;
  wire[6:0] pcr_io_status_zero;
  wire pcr_io_status_er;
  wire pcr_io_status_vm;
  wire pcr_io_status_s64;
  wire pcr_io_status_u64;
  wire pcr_io_status_ef;
  wire pcr_io_status_pei;
  wire pcr_io_status_ei;
  wire pcr_io_status_ps;
  wire pcr_io_status_s;
  wire[31:0] pcr_io_ptbr;
  wire[43:0] pcr_io_evec;
  wire pcr_io_fatc;
  wire pcr_io_replay;
  wire[63:0] pcr_io_time;
  wire[2:0] pcr_io_fcsr_rm;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_kill = {1{$random}};
    mem_reg_kill = {1{$random}};
    R10 = {2{$random}};
    R11 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T18[initvar] = {2{$random}};
    wb_reg_wdata = {2{$random}};
    mem_reg_wdata = {2{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R93 = {2{$random}};
    R94 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    R143 = {1{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T7 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T6 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign T5 = io_ctrl_killd ^ 1'h1;
  assign T6 = ex_reg_kill ^ 1'h1;
  assign T7 = mem_reg_kill ^ 1'h1;
  assign T8 = wb_reg_inst;
  assign T9 = R10;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T82 : T12;
  assign T12 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T13 = T77 ? io_ctrl_bypass_src_1 : T14;
  assign T14 = T76 ? T15 : ex_reg_rs_lsb_1;
  assign T15 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T16;
  assign T16 = T74 ? wb_wdata : T17;
  assign T17 = T18[T26];
  assign T20 = T23 & T21;
  assign T21 = T22 < 5'h1f;
  assign T22 = T25[3'h4:1'h0];
  assign T23 = wb_wen & T24;
  assign T24 = wb_waddr != 5'h0;
  assign wb_waddr = io_ctrl_ll_wen ? io_ctrl_ll_waddr : io_ctrl_wb_waddr;
  assign wb_wen = io_ctrl_ll_wen | io_ctrl_wb_wen;
  assign T25 = ~ wb_waddr;
  assign T26 = ~ T27;
  assign T27 = io_imem_resp_bits_data_0[5'h18:5'h14];
  assign wb_wdata = T28;
  assign T28 = T71 ? io_dmem_resp_bits_data_subword : T29;
  assign T29 = io_ctrl_ll_wen ? ll_wdata : T30;
  assign T30 = T70 ? pcr_io_rw_rdata : wb_reg_wdata;
  assign T31 = T7 ? T32 : wb_reg_wdata;
  assign T32 = T69 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = io_ctrl_mem_ctrl_jalr ? T281 : mem_reg_wdata;
  assign T33 = T6 ? alu_io_out : mem_reg_wdata;
  assign T281 = {T288, mem_br_target};
  assign mem_br_target = T282 + T34;
  assign T34 = T35;
  assign T35 = {1'h0, mem_reg_pc};
  assign T36 = T6 ? ex_reg_pc : mem_reg_pc;
  assign T37 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T282 = {T286, T38};
  assign T38 = T68 ? T283 : T39;
  assign T39 = io_ctrl_mem_ctrl_jal ? T40 : 22'h4;
  assign T40 = T41;
  assign T41 = {T49, T42};
  assign T42 = {T45, T43};
  assign T43 = {T44, 1'h0};
  assign T44 = mem_reg_inst[5'h18:5'h15];
  assign T45 = {T47, T46};
  assign T46 = mem_reg_inst[5'h1e:5'h19];
  assign T47 = T48;
  assign T48 = mem_reg_inst[5'h14:5'h14];
  assign T49 = {T53, T50};
  assign T50 = {T53, T51};
  assign T51 = T52;
  assign T52 = mem_reg_inst[5'h13:4'hc];
  assign T53 = T54;
  assign T54 = mem_reg_inst[5'h1f:5'h1f];
  assign T283 = {T284, T55};
  assign T55 = T56;
  assign T56 = {T64, T57};
  assign T57 = {T60, T58};
  assign T58 = {T59, 1'h0};
  assign T59 = mem_reg_inst[4'hb:4'h8];
  assign T60 = {T62, T61};
  assign T61 = mem_reg_inst[5'h1e:5'h19];
  assign T62 = T63;
  assign T63 = mem_reg_inst[3'h7:3'h7];
  assign T64 = {T66, T65};
  assign T65 = {T66, T66};
  assign T66 = T67;
  assign T67 = mem_reg_inst[5'h1f:5'h1f];
  assign T284 = T285 ? 7'h7f : 7'h0;
  assign T285 = T55[4'he:4'he];
  assign T68 = io_ctrl_mem_ctrl_branch & io_ctrl_mem_br_taken;
  assign T286 = T287 ? 23'h7fffff : 23'h0;
  assign T287 = T38[5'h15:5'h15];
  assign T288 = T289 ? 19'h7ffff : 19'h0;
  assign T289 = mem_br_target[6'h2c:6'h2c];
  assign T69 = io_ctrl_mem_ctrl_fp & io_ctrl_mem_ctrl_wxd;
  assign T70 = io_ctrl_csr != 3'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign T71 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_xpu = T72 ^ 1'h1;
  assign T72 = T73;
  assign T73 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T74 = T23 & T75;
  assign T75 = wb_waddr == T27;
  assign T76 = T5 & io_ctrl_ren_1;
  assign T77 = T5 & io_ctrl_bypass_1;
  assign T78 = T80 ? T79 : ex_reg_rs_msb_1;
  assign T79 = id_rs_1 >> 2'h2;
  assign T80 = T76 & T81;
  assign T81 = io_ctrl_bypass_1 ^ 1'h1;
  assign T82 = T88 ? T86 : T83;
  assign T83 = T84 ? bypass_1 : T290;
  assign T290 = {63'h0, bypass_0};
  assign bypass_0 = 1'h0;
  assign bypass_1 = mem_reg_wdata;
  assign T84 = T85[1'h0:1'h0];
  assign T85 = ex_reg_rs_lsb_1;
  assign T86 = T87 ? bypass_3 : bypass_2;
  assign bypass_2 = wb_reg_wdata;
  assign bypass_3 = io_dmem_resp_bits_data;
  assign T87 = T85[1'h0:1'h0];
  assign T88 = T85[1'h1:1'h1];
  assign T89 = T5 ? io_ctrl_bypass_1 : ex_reg_rs_bypass_1;
  assign T90 = T91;
  assign T91 = wb_reg_inst[5'h18:5'h14];
  assign T92 = R93;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T111 : T95;
  assign T95 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T96 = T106 ? io_ctrl_bypass_src_0 : T97;
  assign T97 = T105 ? T98 : ex_reg_rs_lsb_0;
  assign T98 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T99;
  assign T99 = T103 ? wb_wdata : T100;
  assign T100 = T18[T101];
  assign T101 = ~ T102;
  assign T102 = io_imem_resp_bits_data_0[5'h13:4'hf];
  assign T103 = T23 & T104;
  assign T104 = wb_waddr == T102;
  assign T105 = T5 & io_ctrl_ren_0;
  assign T106 = T5 & io_ctrl_bypass_0;
  assign T107 = T109 ? T108 : ex_reg_rs_msb_0;
  assign T108 = id_rs_0 >> 2'h2;
  assign T109 = T105 & T110;
  assign T110 = io_ctrl_bypass_0 ^ 1'h1;
  assign T111 = T117 ? T115 : T112;
  assign T112 = T113 ? bypass_1 : T291;
  assign T291 = {63'h0, bypass_0};
  assign T113 = T114[1'h0:1'h0];
  assign T114 = ex_reg_rs_lsb_0;
  assign T115 = T116 ? bypass_3 : bypass_2;
  assign T116 = T114[1'h0:1'h0];
  assign T117 = T114[1'h1:1'h1];
  assign T118 = T5 ? io_ctrl_bypass_0 : ex_reg_rs_bypass_0;
  assign T119 = T120;
  assign T120 = wb_reg_inst[5'h13:4'hf];
  assign T121 = wb_wen;
  assign T122 = wb_wdata;
  assign T123 = T124;
  assign T124 = wb_wen ? wb_waddr : 5'h0;
  assign T125 = wb_reg_pc;
  assign T126 = T7 ? mem_reg_pc : wb_reg_pc;
  assign T127 = io_ctrl_retire;
  assign T128 = T129;
  assign T129 = pcr_io_time[6'h20:1'h0];
  assign T130 = io_host_id;
  assign T132 = T138 ? T137 : T133;
  assign T133 = T136 ? T134 : wb_reg_wdata;
  assign T134 = pcr_io_rw_rdata & T135;
  assign T135 = ~ wb_reg_wdata;
  assign T136 = io_ctrl_csr == 3'h3;
  assign T137 = pcr_io_rw_rdata | wb_reg_wdata;
  assign T138 = io_ctrl_csr == 3'h2;
  assign T292 = io_ctrl_csr[1'h1:1'h0];
  assign T139 = wb_reg_inst[5'h1f:5'h14];
  assign T140 = T141 ? 1'h0 : io_ctrl_ll_ready;
  assign T141 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T142 = io_ctrl_killm & R143;
  assign T144 = div_io_req_ready & T145;
  assign T145 = io_ctrl_ex_valid & io_ctrl_ex_ctrl_div;
  assign ex_op1 = T150 ? T149 : T293;
  assign T293 = {T294, T146};
  assign T146 = T148 ? T147 : 44'h0;
  assign T147 = ex_reg_pc;
  assign T148 = io_ctrl_ex_ctrl_sel_alu1 == 2'h2;
  assign T294 = T295 ? 20'hfffff : 20'h0;
  assign T295 = T146[6'h2b:6'h2b];
  assign T149 = ex_rs_0;
  assign T150 = io_ctrl_ex_ctrl_sel_alu1 == 2'h1;
  assign T151 = ex_op2;
  assign ex_op2 = T212 ? T211 : T296;
  assign T296 = {T302, T152};
  assign T152 = T210 ? ex_imm : T297;
  assign T297 = {T298, T153};
  assign T153 = T154 ? 4'h4 : 4'h0;
  assign T154 = io_ctrl_ex_ctrl_sel_alu2 == 2'h1;
  assign T298 = T299 ? 28'hfffffff : 28'h0;
  assign T299 = T153[2'h3:2'h3];
  assign ex_imm = T155;
  assign T155 = {T198, T156};
  assign T156 = {T178, T157};
  assign T157 = {T167, T158};
  assign T158 = T166 ? T165 : T159;
  assign T159 = T164 ? T163 : T160;
  assign T160 = T162 ? T161 : 1'h0;
  assign T161 = ex_reg_inst[4'hf:4'hf];
  assign T162 = io_ctrl_ex_ctrl_sel_imm == 3'h5;
  assign T163 = ex_reg_inst[5'h14:5'h14];
  assign T164 = io_ctrl_ex_ctrl_sel_imm == 3'h4;
  assign T165 = ex_reg_inst[3'h7:3'h7];
  assign T166 = io_ctrl_ex_ctrl_sel_imm == 3'h0;
  assign T167 = T177 ? 4'h0 : T168;
  assign T168 = T174 ? T173 : T169;
  assign T169 = T172 ? T171 : T170;
  assign T170 = ex_reg_inst[5'h18:5'h15];
  assign T171 = ex_reg_inst[5'h13:5'h10];
  assign T172 = io_ctrl_ex_ctrl_sel_imm == 3'h5;
  assign T173 = ex_reg_inst[4'hb:4'h8];
  assign T174 = T176 | T175;
  assign T175 = io_ctrl_ex_ctrl_sel_imm == 3'h1;
  assign T176 = io_ctrl_ex_ctrl_sel_imm == 3'h0;
  assign T177 = io_ctrl_ex_ctrl_sel_imm == 3'h2;
  assign T178 = {T184, T179};
  assign T179 = T181 ? 6'h0 : T180;
  assign T180 = ex_reg_inst[5'h1e:5'h19];
  assign T181 = T183 | T182;
  assign T182 = io_ctrl_ex_ctrl_sel_imm == 3'h5;
  assign T183 = io_ctrl_ex_ctrl_sel_imm == 3'h2;
  assign T184 = T195 ? 1'h0 : T185;
  assign T185 = T194 ? T192 : T186;
  assign T186 = T191 ? T189 : T187;
  assign T187 = T188;
  assign T188 = ex_reg_inst[5'h1f:5'h1f];
  assign T189 = T190;
  assign T190 = ex_reg_inst[3'h7:3'h7];
  assign T191 = io_ctrl_ex_ctrl_sel_imm == 3'h1;
  assign T192 = T193;
  assign T193 = ex_reg_inst[5'h14:5'h14];
  assign T194 = io_ctrl_ex_ctrl_sel_imm == 3'h3;
  assign T195 = T197 | T196;
  assign T196 = io_ctrl_ex_ctrl_sel_imm == 3'h5;
  assign T197 = io_ctrl_ex_ctrl_sel_imm == 3'h2;
  assign T198 = {T187, T199};
  assign T199 = {T206, T200};
  assign T200 = T203 ? T300 : T201;
  assign T201 = T202;
  assign T202 = ex_reg_inst[5'h13:4'hc];
  assign T300 = T187 ? 8'hff : 8'h0;
  assign T203 = T205 & T204;
  assign T204 = io_ctrl_ex_ctrl_sel_imm != 3'h3;
  assign T205 = io_ctrl_ex_ctrl_sel_imm != 3'h2;
  assign T206 = T209 ? T207 : T301;
  assign T301 = T187 ? 11'h7ff : 11'h0;
  assign T207 = T208;
  assign T208 = ex_reg_inst[5'h1e:5'h14];
  assign T209 = io_ctrl_ex_ctrl_sel_imm == 3'h2;
  assign T210 = io_ctrl_ex_ctrl_sel_alu2 == 2'h3;
  assign T302 = T303 ? 32'hffffffff : 32'h0;
  assign T303 = T152[5'h1f:5'h1f];
  assign T211 = ex_rs_1;
  assign T212 = io_ctrl_ex_ctrl_sel_alu2 == 2'h2;
//  assign io_rocc_exception = {1{$random}};
//  assign io_rocc_pptw_sret = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_s = {1{$random}};
//  assign io_rocc_pptw_status_ps = {1{$random}};
//  assign io_rocc_pptw_status_ei = {1{$random}};
//  assign io_rocc_pptw_status_pei = {1{$random}};
//  assign io_rocc_pptw_status_ef = {1{$random}};
//  assign io_rocc_pptw_status_u64 = {1{$random}};
//  assign io_rocc_pptw_status_s64 = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_er = {1{$random}};
//  assign io_rocc_pptw_status_zero = {1{$random}};
//  assign io_rocc_pptw_status_im = {1{$random}};
//  assign io_rocc_pptw_status_ip = {1{$random}};
//  assign io_rocc_pptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_pptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_sret = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_s = {1{$random}};
//  assign io_rocc_dptw_status_ps = {1{$random}};
//  assign io_rocc_dptw_status_ei = {1{$random}};
//  assign io_rocc_dptw_status_pei = {1{$random}};
//  assign io_rocc_dptw_status_ef = {1{$random}};
//  assign io_rocc_dptw_status_u64 = {1{$random}};
//  assign io_rocc_dptw_status_s64 = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_er = {1{$random}};
//  assign io_rocc_dptw_status_zero = {1{$random}};
//  assign io_rocc_dptw_status_im = {1{$random}};
//  assign io_rocc_dptw_status_ip = {1{$random}};
//  assign io_rocc_dptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_dptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_sret = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_s = {1{$random}};
//  assign io_rocc_iptw_status_ps = {1{$random}};
//  assign io_rocc_iptw_status_ei = {1{$random}};
//  assign io_rocc_iptw_status_pei = {1{$random}};
//  assign io_rocc_iptw_status_ef = {1{$random}};
//  assign io_rocc_iptw_status_u64 = {1{$random}};
//  assign io_rocc_iptw_status_s64 = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_er = {1{$random}};
//  assign io_rocc_iptw_status_zero = {1{$random}};
//  assign io_rocc_iptw_status_im = {1{$random}};
//  assign io_rocc_iptw_status_ip = {1{$random}};
//  assign io_rocc_iptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_iptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_release_ready = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_p_type = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_addr = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_probe_valid = {1{$random}};
//  assign io_rocc_dmem_finish_ready = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_dmem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_grant_valid = {1{$random}};
//  assign io_rocc_dmem_acquire_ready = {1{$random}};
//  assign io_rocc_imem_finish_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_imem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_imem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
//  assign io_rocc_s = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_ptw_req_bits = {1{$random}};
//  assign io_rocc_mem_ptw_req_valid = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_data_subword = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T213 = T218 ? mem_reg_rs2 : wb_reg_rs2;
  assign T214 = T215 ? ex_rs_1 : mem_reg_rs2;
  assign T215 = T6 & T216;
  assign T216 = io_ctrl_ex_ctrl_rxs2 & T217;
  assign T217 = io_ctrl_ex_ctrl_mem | io_ctrl_ex_ctrl_rocc;
  assign T218 = T7 & io_ctrl_mem_ctrl_rocc;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_inst_opcode = T219;
  assign T219 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T220;
  assign T220 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T221;
  assign T221 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T222;
  assign T222 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T223;
  assign T223 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T224;
  assign T224 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T225;
  assign T225 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T226;
  assign T226 = wb_reg_inst[5'h1f:5'h19];
//  assign io_rocc_cmd_valid = {1{$random}};
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = T304;
  assign T304 = dmem_resp_waddr[3'h4:1'h0];
  assign dmem_resp_waddr = T227 >> 1'h1;
  assign T227 = io_dmem_resp_bits_tag;
  assign io_fpu_dmem_resp_type = T305;
  assign T305 = io_dmem_resp_bits_typ[2'h2:1'h0];
  assign io_fpu_dmem_resp_val = T228;
  assign T228 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T229;
  assign T229 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = pcr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
//  assign io_imem_invalidate = {1{$random}};
//  assign io_imem_ptw_sret = {1{$random}};
//  assign io_imem_ptw_invalidate = {1{$random}};
//  assign io_imem_ptw_status_s = {1{$random}};
//  assign io_imem_ptw_status_ps = {1{$random}};
//  assign io_imem_ptw_status_ei = {1{$random}};
//  assign io_imem_ptw_status_pei = {1{$random}};
//  assign io_imem_ptw_status_ef = {1{$random}};
//  assign io_imem_ptw_status_u64 = {1{$random}};
//  assign io_imem_ptw_status_s64 = {1{$random}};
//  assign io_imem_ptw_status_vm = {1{$random}};
//  assign io_imem_ptw_status_er = {1{$random}};
//  assign io_imem_ptw_status_zero = {1{$random}};
//  assign io_imem_ptw_status_im = {1{$random}};
//  assign io_imem_ptw_status_ip = {1{$random}};
//  assign io_imem_ptw_resp_bits_perm = {1{$random}};
//  assign io_imem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_imem_ptw_resp_bits_error = {1{$random}};
//  assign io_imem_ptw_resp_valid = {1{$random}};
//  assign io_imem_ptw_req_ready = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_bht_value = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_bht_history = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_entry = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_target = {2{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_bridx = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_mask = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_bits_taken = {1{$random}};
//  assign io_imem_ras_update_bits_prediction_valid = {1{$random}};
  assign io_imem_ras_update_bits_returnAddr = T306;
  assign T306 = mem_int_wdata[6'h2a:1'h0];
//  assign io_imem_ras_update_bits_isReturn = {1{$random}};
//  assign io_imem_ras_update_bits_isCall = {1{$random}};
//  assign io_imem_ras_update_valid = {1{$random}};
//  assign io_imem_bht_update_bits_mispredict = {1{$random}};
//  assign io_imem_bht_update_bits_taken = {1{$random}};
  assign io_imem_bht_update_bits_pc = T307;
  assign T307 = mem_reg_pc[6'h2a:1'h0];
//  assign io_imem_bht_update_bits_prediction_bits_bht_value = {1{$random}};
//  assign io_imem_bht_update_bits_prediction_bits_bht_history = {1{$random}};
//  assign io_imem_bht_update_bits_prediction_bits_entry = {1{$random}};
//  assign io_imem_bht_update_bits_prediction_bits_target = {2{$random}};
//  assign io_imem_bht_update_bits_prediction_bits_bridx = {1{$random}};
//  assign io_imem_bht_update_bits_prediction_bits_mask = {1{$random}};
//  assign io_imem_bht_update_bits_prediction_bits_taken = {1{$random}};
//  assign io_imem_bht_update_bits_prediction_valid = {1{$random}};
//  assign io_imem_bht_update_valid = {1{$random}};
  assign io_imem_btb_update_bits_br_pc = T308;
  assign T308 = mem_reg_pc[6'h2a:1'h0];
//  assign io_imem_btb_update_bits_isReturn = {1{$random}};
//  assign io_imem_btb_update_bits_isJump = {1{$random}};
//  assign io_imem_btb_update_bits_taken = {1{$random}};
  assign io_imem_btb_update_bits_target = T309;
  assign T309 = io_imem_req_bits_pc[6'h2a:1'h0];
  assign io_imem_btb_update_bits_pc = T310;
  assign T310 = mem_reg_pc[6'h2a:1'h0];
//  assign io_imem_btb_update_bits_prediction_bits_bht_value = {1{$random}};
//  assign io_imem_btb_update_bits_prediction_bits_bht_history = {1{$random}};
//  assign io_imem_btb_update_bits_prediction_bits_entry = {1{$random}};
//  assign io_imem_btb_update_bits_prediction_bits_target = {2{$random}};
//  assign io_imem_btb_update_bits_prediction_bits_bridx = {1{$random}};
//  assign io_imem_btb_update_bits_prediction_bits_mask = {1{$random}};
//  assign io_imem_btb_update_bits_prediction_bits_taken = {1{$random}};
//  assign io_imem_btb_update_bits_prediction_valid = {1{$random}};
//  assign io_imem_btb_update_valid = {1{$random}};
//  assign io_imem_resp_ready = {1{$random}};
  assign io_imem_req_bits_pc = T311;
  assign T311 = T230[6'h2b:1'h0];
  assign T230 = T231;
  assign T231 = T249 ? mem_npc : T312;
  assign T312 = {1'h0, T232};
  assign T232 = T233 ? pcr_io_evec : wb_reg_pc;
  assign T233 = io_ctrl_sel_pc == 3'h3;
  assign mem_npc = io_ctrl_mem_ctrl_jalr ? T313 : mem_br_target;
  assign T313 = {1'h0, T234};
  assign T234 = {T236, T235};
  assign T235 = mem_reg_wdata[6'h2a:1'h0];
  assign T236 = T246 ? T245 : T237;
  assign T237 = T241 ? T240 : T238;
  assign T238 = T239[1'h0:1'h0];
  assign T239 = mem_reg_wdata[6'h2b:6'h2a];
  assign T240 = T239 == 2'h3;
  assign T241 = T244 | T242;
  assign T242 = T243 == 22'h3ffffe;
  assign T243 = mem_reg_wdata >> 6'h2a;
  assign T244 = T243 == 22'h3fffff;
  assign T245 = T239 != 2'h0;
  assign T246 = T248 | T247;
  assign T247 = T243 == 22'h1;
  assign T248 = T243 == 22'h0;
  assign T249 = io_ctrl_sel_pc == 3'h1;
//  assign io_imem_req_valid = {1{$random}};
  assign io_ptw_status_s = pcr_io_status_s;
  assign io_ptw_status_ps = pcr_io_status_ps;
  assign io_ptw_status_ei = pcr_io_status_ei;
  assign io_ptw_status_pei = pcr_io_status_pei;
  assign io_ptw_status_ef = pcr_io_status_ef;
  assign io_ptw_status_u64 = pcr_io_status_u64;
  assign io_ptw_status_s64 = pcr_io_status_s64;
  assign io_ptw_status_vm = pcr_io_status_vm;
  assign io_ptw_status_er = pcr_io_status_er;
  assign io_ptw_status_zero = pcr_io_status_zero;
  assign io_ptw_status_im = pcr_io_status_im;
  assign io_ptw_status_ip = pcr_io_status_ip;
  assign io_ptw_sret = io_ctrl_sret;
  assign io_ptw_invalidate = pcr_io_fatc;
  assign io_ptw_ptbr = pcr_io_ptbr;
//  assign io_dmem_ptw_sret = {1{$random}};
//  assign io_dmem_ptw_invalidate = {1{$random}};
//  assign io_dmem_ptw_status_s = {1{$random}};
//  assign io_dmem_ptw_status_ps = {1{$random}};
//  assign io_dmem_ptw_status_ei = {1{$random}};
//  assign io_dmem_ptw_status_pei = {1{$random}};
//  assign io_dmem_ptw_status_ef = {1{$random}};
//  assign io_dmem_ptw_status_u64 = {1{$random}};
//  assign io_dmem_ptw_status_s64 = {1{$random}};
//  assign io_dmem_ptw_status_vm = {1{$random}};
//  assign io_dmem_ptw_status_er = {1{$random}};
//  assign io_dmem_ptw_status_zero = {1{$random}};
//  assign io_dmem_ptw_status_im = {1{$random}};
//  assign io_dmem_ptw_status_ip = {1{$random}};
//  assign io_dmem_ptw_resp_bits_perm = {1{$random}};
//  assign io_dmem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_dmem_ptw_resp_bits_error = {1{$random}};
//  assign io_dmem_ptw_resp_valid = {1{$random}};
//  assign io_dmem_ptw_req_ready = {1{$random}};
  assign io_dmem_req_bits_data = T250;
  assign T250 = io_ctrl_mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
//  assign io_dmem_req_bits_cmd = {1{$random}};
  assign io_dmem_req_bits_tag = T314;
  assign T314 = {2'h0, T251};
  assign T251 = {io_ctrl_ex_waddr, io_ctrl_ex_ctrl_fp};
  assign io_dmem_req_bits_addr = T252;
  assign T252 = T253;
  assign T253 = {T255, T254};
  assign T254 = alu_io_adder_out[6'h2a:1'h0];
  assign T255 = T265 ? T264 : T256;
  assign T256 = T260 ? T259 : T257;
  assign T257 = T258[1'h0:1'h0];
  assign T258 = alu_io_adder_out[6'h2b:6'h2a];
  assign T259 = T258 == 2'h3;
  assign T260 = T263 | T261;
  assign T261 = T262 == 22'h3ffffe;
  assign T262 = ex_rs_0 >> 6'h2a;
  assign T263 = T262 == 22'h3fffff;
  assign T264 = T258 != 2'h0;
  assign T265 = T267 | T266;
  assign T266 = T262 == 22'h1;
  assign T267 = T262 == 22'h0;
//  assign io_dmem_req_bits_phys = {1{$random}};
//  assign io_dmem_req_bits_typ = {1{$random}};
//  assign io_dmem_req_bits_kill = {1{$random}};
//  assign io_dmem_req_valid = {1{$random}};
  assign io_ctrl_csr_replay = pcr_io_replay;
  assign io_ctrl_fp_sboard_clra = T315;
  assign T315 = dmem_resp_waddr[3'h4:1'h0];
  assign io_ctrl_fp_sboard_clr = T268;
  assign T268 = dmem_resp_replay & dmem_resp_fpu;
  assign io_ctrl_status_s = pcr_io_status_s;
  assign io_ctrl_status_ps = pcr_io_status_ps;
  assign io_ctrl_status_ei = pcr_io_status_ei;
  assign io_ctrl_status_pei = pcr_io_status_pei;
  assign io_ctrl_status_ef = pcr_io_status_ef;
  assign io_ctrl_status_u64 = pcr_io_status_u64;
  assign io_ctrl_status_s64 = pcr_io_status_s64;
  assign io_ctrl_status_vm = pcr_io_status_vm;
  assign io_ctrl_status_er = pcr_io_status_er;
  assign io_ctrl_status_zero = pcr_io_status_zero;
  assign io_ctrl_status_im = pcr_io_status_im;
  assign io_ctrl_status_ip = pcr_io_status_ip;
  assign io_ctrl_wb_waddr = T269;
  assign T269 = wb_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_waddr = T270;
  assign T270 = mem_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_rs1_ra = T271;
  assign T271 = T272 == 5'h1;
  assign T272 = mem_reg_inst[5'h13:4'hf];
  assign io_ctrl_ex_waddr = T273;
  assign T273 = ex_reg_inst[4'hb:3'h7];
  assign io_ctrl_ll_waddr = T316;
  assign T316 = T274[3'h4:1'h0];
  assign T274 = T141 ? dmem_resp_waddr : T317;
  assign T317 = {2'h0, div_io_resp_bits_tag};
  assign io_ctrl_ll_wen = T275;
  assign T275 = T141 ? 1'h1 : T276;
  assign T276 = T140 & div_io_resp_valid;
  assign io_ctrl_div_mul_rdy = div_io_req_ready;
  assign io_ctrl_mem_misprediction = T277;
  assign T277 = T279 | T278;
  assign T278 = io_ctrl_ex_valid ^ 1'h1;
  assign T279 = mem_npc != T318;
  assign T318 = {1'h0, ex_reg_pc};
  assign io_ctrl_mem_br_taken = T280;
  assign T280 = mem_reg_wdata[1'h0:1'h0];
  assign io_ctrl_inst = io_imem_resp_bits_data_0;
  assign io_host_debug_stats_pcr = pcr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = pcr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = pcr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = pcr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = pcr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = pcr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = pcr_io_host_pcr_req_ready;
  ALU alu(
       .io_dw( io_ctrl_ex_ctrl_alu_dw ),
       .io_fn( io_ctrl_ex_ctrl_alu_fn ),
       .io_in2( T151 ),
       .io_in1( ex_op1 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( T145 ),
       .io_req_bits_fn( io_ctrl_ex_ctrl_alu_fn ),
       .io_req_bits_dw( io_ctrl_ex_ctrl_alu_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( io_ctrl_ex_waddr ),
       .io_kill( T142 ),
       .io_resp_ready( T140 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );
  CSRFile pcr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( pcr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( pcr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( pcr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( pcr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( pcr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( pcr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( pcr_io_host_debug_stats_pcr ),
       .io_rw_addr( T139 ),
       .io_rw_cmd( T292 ),
       .io_rw_rdata( pcr_io_rw_rdata ),
       .io_rw_wdata( T132 ),
       .io_status_ip( pcr_io_status_ip ),
       .io_status_im( pcr_io_status_im ),
       .io_status_zero( pcr_io_status_zero ),
       .io_status_er( pcr_io_status_er ),
       .io_status_vm( pcr_io_status_vm ),
       .io_status_s64( pcr_io_status_s64 ),
       .io_status_u64( pcr_io_status_u64 ),
       .io_status_ef( pcr_io_status_ef ),
       .io_status_pei( pcr_io_status_pei ),
       .io_status_ei( pcr_io_status_ei ),
       .io_status_ps( pcr_io_status_ps ),
       .io_status_s( pcr_io_status_s ),
       .io_ptbr( pcr_io_ptbr ),
       .io_evec( pcr_io_evec ),
       .io_exception( io_ctrl_exception ),
       .io_retire( io_ctrl_retire ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( io_ctrl_cause ),
       .io_badvaddr_wen( io_ctrl_badvaddr_wen ),
       .io_pc( wb_reg_pc ),
       .io_sret( io_ctrl_sret ),
       .io_fatc( pcr_io_fatc ),
       .io_replay( pcr_io_replay ),
       .io_time( pcr_io_time ),
       .io_fcsr_rm( pcr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_manager_xact_id( io_rocc_imem_finish_bits_payload_manager_xact_id ),
       //.io_rocc_dmem_acquire_ready(  )
       .io_rocc_dmem_acquire_valid( io_rocc_dmem_acquire_valid ),
       .io_rocc_dmem_acquire_bits_header_src( io_rocc_dmem_acquire_bits_header_src ),
       .io_rocc_dmem_acquire_bits_header_dst( io_rocc_dmem_acquire_bits_header_dst ),
       .io_rocc_dmem_acquire_bits_payload_addr( io_rocc_dmem_acquire_bits_payload_addr ),
       .io_rocc_dmem_acquire_bits_payload_client_xact_id( io_rocc_dmem_acquire_bits_payload_client_xact_id ),
       .io_rocc_dmem_acquire_bits_payload_data( io_rocc_dmem_acquire_bits_payload_data ),
       .io_rocc_dmem_acquire_bits_payload_uncached( io_rocc_dmem_acquire_bits_payload_uncached ),
       .io_rocc_dmem_acquire_bits_payload_a_type( io_rocc_dmem_acquire_bits_payload_a_type ),
       .io_rocc_dmem_acquire_bits_payload_subblock( io_rocc_dmem_acquire_bits_payload_subblock ),
       .io_rocc_dmem_grant_ready( io_rocc_dmem_grant_ready ),
       //.io_rocc_dmem_grant_valid(  )
       //.io_rocc_dmem_grant_bits_header_src(  )
       //.io_rocc_dmem_grant_bits_header_dst(  )
       //.io_rocc_dmem_grant_bits_payload_data(  )
       //.io_rocc_dmem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_uncached(  )
       //.io_rocc_dmem_grant_bits_payload_g_type(  )
       //.io_rocc_dmem_finish_ready(  )
       .io_rocc_dmem_finish_valid( io_rocc_dmem_finish_valid ),
       .io_rocc_dmem_finish_bits_header_src( io_rocc_dmem_finish_bits_header_src ),
       .io_rocc_dmem_finish_bits_header_dst( io_rocc_dmem_finish_bits_header_dst ),
       .io_rocc_dmem_finish_bits_payload_manager_xact_id( io_rocc_dmem_finish_bits_payload_manager_xact_id ),
       .io_rocc_dmem_probe_ready( io_rocc_dmem_probe_ready ),
       //.io_rocc_dmem_probe_valid(  )
       //.io_rocc_dmem_probe_bits_header_src(  )
       //.io_rocc_dmem_probe_bits_header_dst(  )
       //.io_rocc_dmem_probe_bits_payload_addr(  )
       //.io_rocc_dmem_probe_bits_payload_p_type(  )
       //.io_rocc_dmem_release_ready(  )
       .io_rocc_dmem_release_valid( io_rocc_dmem_release_valid ),
       .io_rocc_dmem_release_bits_header_src( io_rocc_dmem_release_bits_header_src ),
       .io_rocc_dmem_release_bits_header_dst( io_rocc_dmem_release_bits_header_dst ),
       .io_rocc_dmem_release_bits_payload_addr( io_rocc_dmem_release_bits_payload_addr ),
       .io_rocc_dmem_release_bits_payload_client_xact_id( io_rocc_dmem_release_bits_payload_client_xact_id ),
       .io_rocc_dmem_release_bits_payload_data( io_rocc_dmem_release_bits_payload_data ),
       .io_rocc_dmem_release_bits_payload_r_type( io_rocc_dmem_release_bits_payload_r_type ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );

  always @(posedge clk) begin
    if(T7) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T6) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data_0;
    end
    ex_reg_kill <= io_ctrl_killd;
    mem_reg_kill <= ex_reg_kill;
    R10 <= R11;
    if(ex_reg_rs_bypass_1) begin
      R11 <= T82;
    end else begin
      R11 <= T12;
    end
    if(T77) begin
      ex_reg_rs_lsb_1 <= io_ctrl_bypass_src_1;
    end else if(T76) begin
      ex_reg_rs_lsb_1 <= T15;
    end
    if (T20)
      T18[T25] <= wb_wdata;
    if(T7) begin
      wb_reg_wdata <= T32;
    end
    if(T6) begin
      mem_reg_wdata <= alu_io_out;
    end
    if(T6) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T80) begin
      ex_reg_rs_msb_1 <= T79;
    end
    if(T5) begin
      ex_reg_rs_bypass_1 <= io_ctrl_bypass_1;
    end
    R93 <= R94;
    if(ex_reg_rs_bypass_0) begin
      R94 <= T111;
    end else begin
      R94 <= T95;
    end
    if(T106) begin
      ex_reg_rs_lsb_0 <= io_ctrl_bypass_src_0;
    end else if(T105) begin
      ex_reg_rs_lsb_0 <= T98;
    end
    if(T109) begin
      ex_reg_rs_msb_0 <= T108;
    end
    if(T5) begin
      ex_reg_rs_bypass_0 <= io_ctrl_bypass_0;
    end
    if(T7) begin
      wb_reg_pc <= mem_reg_pc;
    end
    R143 <= T144;
    if(T218) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(T215) begin
      mem_reg_rs2 <= ex_rs_1;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T130, T128, T127, T125, T123, T122, T121, T119, T92, T90, T9, T8, T1);
// synthesis translate_on
`endif
  end
endmodule

module FPUDecoder(
    input [31:0] io_inst,
    output[4:0] io_sigs_cmd,
    output io_sigs_ldst,
    output io_sigs_wen,
    output io_sigs_ren1,
    output io_sigs_ren2,
    output io_sigs_ren3,
    output io_sigs_swap23,
    output io_sigs_single,
    output io_sigs_fromint,
    output io_sigs_toint,
    output io_sigs_fastpipe,
    output io_sigs_fma,
    output io_sigs_round
);

  wire T0;
  wire T1;
  wire[31:0] T2;
  wire T3;
  wire T4;
  wire[31:0] T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  wire T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire T16;
  wire[31:0] T17;
  wire T18;
  wire T19;
  wire[31:0] T20;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire[31:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire T41;
  wire[31:0] T42;
  wire T43;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire[31:0] T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire[31:0] T55;
  wire T56;
  wire T57;
  wire[31:0] T58;
  wire T59;
  wire T60;
  wire[31:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[31:0] T65;
  wire T66;
  wire T67;
  wire[31:0] T68;
  wire T69;
  wire T70;
  wire[31:0] T71;
  wire T72;
  wire T73;
  wire[31:0] T74;
  wire T75;
  wire T76;
  wire[31:0] T77;
  wire T78;
  wire T79;
  wire[31:0] T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[31:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire[31:0] T114;
  wire[4:0] T115;
  wire[3:0] T116;
  wire[2:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire[31:0] T121;
  wire T122;
  wire[31:0] T123;
  wire T124;
  wire T125;
  wire[31:0] T126;
  wire T127;
  wire[31:0] T128;
  wire T129;
  wire T130;
  wire[31:0] T131;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire T135;
  wire[31:0] T136;
  wire T137;
  wire[31:0] T138;


  assign io_sigs_round = T0;
  assign T0 = T3 | T1;
  assign T1 = T2 == 32'he0000053;
  assign T2 = io_inst & 32'hedf0707f;
  assign T3 = T6 | T4;
  assign T4 = T5 == 32'he0000053;
  assign T5 = io_inst & 32'hfdf0607f;
  assign T6 = T9 | T7;
  assign T7 = T8 == 32'hc0000053;
  assign T8 = io_inst & 32'hedc0007f;
  assign T9 = T12 | T10;
  assign T10 = T11 == 32'h42000053;
  assign T11 = io_inst & 32'h7ff0007f;
  assign T12 = T15 | T13;
  assign T13 = T14 == 32'h40100053;
  assign T14 = io_inst & 32'h7ff0007f;
  assign T15 = T18 | T16;
  assign T16 = T17 == 32'h53;
  assign T17 = io_inst & 32'hec00007f;
  assign T18 = T21 | T19;
  assign T19 = T20 == 32'h53;
  assign T20 = io_inst & 32'hf400007f;
  assign T21 = T22 == 32'h43;
  assign T22 = io_inst & 32'h4000073;
  assign io_sigs_fma = T23;
  assign T23 = T24 | T16;
  assign T24 = T21 | T19;
  assign io_sigs_fastpipe = T25;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h42000053;
  assign T27 = io_inst & 32'hfff0007f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h40100053;
  assign T30 = io_inst & 32'hfff0007f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h20000053;
  assign T33 = io_inst & 32'hf400607f;
  assign T34 = T35 == 32'h20000053;
  assign T35 = io_inst & 32'hfc00507f;
  assign io_sigs_toint = T36;
  assign T36 = T37 | T4;
  assign T37 = T40 | T38;
  assign T38 = T39 == 32'hc0000053;
  assign T39 = io_inst & 32'hfdc0007f;
  assign T40 = T43 | T41;
  assign T41 = T42 == 32'ha0000053;
  assign T42 = io_inst & 32'hfc00507f;
  assign T43 = T46 | T44;
  assign T44 = T45 == 32'ha0000053;
  assign T45 = io_inst & 32'hfc00607f;
  assign T46 = T47 == 32'h2027;
  assign T47 = io_inst & 32'h607f;
  assign io_sigs_fromint = T48;
  assign T48 = T51 | T49;
  assign T49 = T50 == 32'hf0000053;
  assign T50 = io_inst & 32'hfdf0707f;
  assign T51 = T52 == 32'hd0000053;
  assign T52 = io_inst & 32'hfdc0007f;
  assign io_sigs_single = T53;
  assign T53 = T56 | T54;
  assign T54 = T55 == 32'he0000053;
  assign T55 = io_inst & 32'heff0707f;
  assign T56 = T59 | T57;
  assign T57 = T58 == 32'he0000053;
  assign T58 = io_inst & 32'hfff0607f;
  assign T59 = T62 | T60;
  assign T60 = T61 == 32'hc0000053;
  assign T61 = io_inst & 32'hefc0007f;
  assign T62 = T63 | T13;
  assign T63 = T66 | T64;
  assign T64 = T65 == 32'h20000053;
  assign T65 = io_inst & 32'h7e00507f;
  assign T66 = T69 | T67;
  assign T67 = T68 == 32'h20000053;
  assign T68 = io_inst & 32'h7e00607f;
  assign T69 = T72 | T70;
  assign T70 = T71 == 32'h20000053;
  assign T71 = io_inst & 32'hf600607f;
  assign T72 = T75 | T73;
  assign T73 = T74 == 32'h2007;
  assign T74 = io_inst & 32'h705f;
  assign T75 = T78 | T76;
  assign T76 = T77 == 32'h53;
  assign T77 = io_inst & 32'hee00007f;
  assign T78 = T81 | T79;
  assign T79 = T80 == 32'h53;
  assign T80 = io_inst & 32'hf600007f;
  assign T81 = T82 == 32'h43;
  assign T82 = io_inst & 32'h6000073;
  assign io_sigs_swap23 = T19;
  assign io_sigs_ren3 = T21;
  assign io_sigs_ren2 = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h20000053;
  assign T85 = io_inst & 32'h7c00507f;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h20000053;
  assign T88 = io_inst & 32'h7c00607f;
  assign T89 = T90 | T32;
  assign T90 = T91 | T46;
  assign T91 = T92 | T16;
  assign T92 = T21 | T19;
  assign io_sigs_ren1 = T93;
  assign T93 = T94 | T4;
  assign T94 = T95 | T38;
  assign T95 = T96 | T10;
  assign T96 = T97 | T13;
  assign T97 = T98 | T84;
  assign T98 = T99 | T87;
  assign T99 = T100 | T32;
  assign T100 = T101 | T16;
  assign T101 = T21 | T19;
  assign io_sigs_wen = T102;
  assign T102 = T103 | T49;
  assign T103 = T104 | T51;
  assign T104 = T105 | T26;
  assign T105 = T106 | T29;
  assign T106 = T107 | T32;
  assign T107 = T108 | T34;
  assign T108 = T111 | T109;
  assign T109 = T110 == 32'h2007;
  assign T110 = io_inst & 32'h607f;
  assign T111 = T112 | T16;
  assign T112 = T21 | T19;
  assign io_sigs_ldst = T113;
  assign T113 = T114 == 32'h2007;
  assign T114 = io_inst & 32'h605f;
  assign io_sigs_cmd = T115;
  assign T115 = {T137, T116};
  assign T116 = {T134, T117};
  assign T117 = {T129, T118};
  assign T118 = {T124, T119};
  assign T119 = T122 | T120;
  assign T120 = T121 == 32'h8000010;
  assign T121 = io_inst & 32'h8000010;
  assign T122 = T123 == 32'h4;
  assign T123 = io_inst & 32'h4;
  assign T124 = T127 | T125;
  assign T125 = T126 == 32'h10000010;
  assign T126 = io_inst & 32'h10000010;
  assign T127 = T128 == 32'h8;
  assign T128 = io_inst & 32'h8;
  assign T129 = T132 | T130;
  assign T130 = T131 == 32'h20000000;
  assign T131 = io_inst & 32'h20000000;
  assign T132 = T133 == 32'h0;
  assign T133 = io_inst & 32'h40;
  assign T134 = T132 | T135;
  assign T135 = T136 == 32'h40000000;
  assign T136 = io_inst & 32'h40000000;
  assign T137 = T138 == 32'h0;
  assign T138 = io_inst & 32'h10;
endmodule

module mulAddSubRecodedFloatN_0(
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[27:0] T4;
  wire[27:0] T529;
  wire[25:0] T5;
  wire[26:0] roundMask;
  wire[26:0] T6;
  wire[24:0] T7;
  wire[24:0] T530;
  wire T8;
  wire[24:0] T9;
  wire[8:0] T10;
  wire T11;
  wire[8:0] T12;
  wire[24:0] T13;
  wire[1024:0] T14;
  wire[9:0] T15;
  wire[9:0] sExpX3_13;
  wire[10:0] sExpX3;
  wire[10:0] T531;
  wire[6:0] estNormDist;
  wire[6:0] T16;
  wire[6:0] estNormNeg_dist;
  wire[6:0] T17;
  wire[6:0] T18;
  wire[6:0] T19;
  wire[6:0] T20;
  wire[6:0] T21;
  wire[6:0] T22;
  wire[6:0] T23;
  wire[6:0] T24;
  wire[6:0] T25;
  wire[6:0] T26;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[6:0] T29;
  wire[6:0] T30;
  wire[6:0] T31;
  wire[6:0] T32;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[6:0] T40;
  wire[6:0] T41;
  wire[6:0] T42;
  wire[6:0] T43;
  wire[6:0] T44;
  wire[6:0] T45;
  wire[6:0] T46;
  wire[6:0] T47;
  wire[6:0] T48;
  wire[6:0] T49;
  wire[6:0] T50;
  wire[6:0] T51;
  wire[6:0] T52;
  wire[6:0] T53;
  wire[6:0] T54;
  wire[6:0] T55;
  wire[6:0] T56;
  wire[6:0] T57;
  wire[6:0] T58;
  wire[6:0] T59;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire T65;
  wire[50:0] T66;
  wire[50:0] T67;
  wire[49:0] T68;
  wire[49:0] T69;
  wire[74:0] sigSum;
  wire[74:0] alignedNegSigC;
  wire[75:0] T70;
  wire T71;
  wire doSubMags;
  wire opSignC;
  wire T72;
  wire T73;
  wire signProd;
  wire T74;
  wire T75;
  wire signB;
  wire signA;
  wire T76;
  wire[23:0] T77;
  wire[23:0] CExtraMask;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[6:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[5:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[3:0] T89;
  wire[7:0] T90;
  wire[23:0] T91;
  wire[128:0] T92;
  wire[6:0] CAlignDist;
  wire[10:0] T93;
  wire[10:0] T94;
  wire[10:0] sNatCAlignDist;
  wire[10:0] T532;
  wire[8:0] expC;
  wire[10:0] sExpAlignedProd;
  wire[10:0] T95;
  wire[10:0] T533;
  wire[8:0] expA;
  wire[10:0] T96;
  wire[7:0] T97;
  wire[8:0] expB;
  wire[2:0] T98;
  wire[2:0] T534;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire CAlignDist_floor;
  wire T103;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T104;
  wire isZeroA;
  wire[2:0] T105;
  wire[7:0] T106;
  wire[7:0] T535;
  wire[3:0] T107;
  wire[7:0] T108;
  wire[7:0] T536;
  wire[5:0] T109;
  wire[7:0] T110;
  wire[7:0] T537;
  wire[6:0] T111;
  wire[15:0] T112;
  wire[15:0] T113;
  wire[15:0] T114;
  wire[14:0] T115;
  wire[15:0] T116;
  wire[15:0] T117;
  wire[15:0] T118;
  wire[13:0] T119;
  wire[15:0] T120;
  wire[15:0] T121;
  wire[15:0] T122;
  wire[11:0] T123;
  wire[15:0] T124;
  wire[15:0] T125;
  wire[15:0] T126;
  wire[7:0] T127;
  wire[15:0] T128;
  wire[15:0] T129;
  wire[15:0] T538;
  wire[7:0] T130;
  wire[15:0] T131;
  wire[15:0] T539;
  wire[11:0] T132;
  wire[15:0] T133;
  wire[15:0] T540;
  wire[13:0] T134;
  wire[15:0] T135;
  wire[15:0] T541;
  wire[14:0] T136;
  wire[23:0] sigC;
  wire[22:0] fractC;
  wire T137;
  wire isZeroC;
  wire[2:0] T138;
  wire[74:0] T139;
  wire[74:0] T140;
  wire[74:0] T141;
  wire[73:0] T142;
  wire[49:0] T143;
  wire[49:0] T542;
  wire[23:0] negSigC;
  wire[23:0] T144;
  wire[74:0] T543;
  wire[48:0] T145;
  wire[47:0] T146;
  wire[23:0] sigB;
  wire[22:0] fractB;
  wire T147;
  wire[23:0] sigA;
  wire[22:0] fractA;
  wire T148;
  wire[50:0] T544;
  wire[49:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire notCDom_signSigSum;
  wire[6:0] CDom_estNormDist;
  wire[6:0] T545;
  wire[4:0] T198;
  wire[6:0] T199;
  wire T200;
  wire CAlignDist_0;
  wire T201;
  wire[9:0] T202;
  wire isCDominant;
  wire T203;
  wire T204;
  wire[9:0] T205;
  wire T206;
  wire[10:0] sExpSum;
  wire[10:0] T546;
  wire[7:0] T207;
  wire[7:0] T208;
  wire[7:0] T209;
  wire[6:0] T210;
  wire[7:0] T211;
  wire[7:0] T212;
  wire[7:0] T213;
  wire[5:0] T214;
  wire[7:0] T215;
  wire[7:0] T216;
  wire[7:0] T217;
  wire[3:0] T218;
  wire[7:0] T219;
  wire[7:0] T220;
  wire[7:0] T547;
  wire[3:0] T221;
  wire[7:0] T222;
  wire[7:0] T548;
  wire[5:0] T223;
  wire[7:0] T224;
  wire[7:0] T549;
  wire[6:0] T225;
  wire[15:0] T226;
  wire[15:0] T227;
  wire[15:0] T228;
  wire[14:0] T229;
  wire[15:0] T230;
  wire[15:0] T231;
  wire[15:0] T232;
  wire[13:0] T233;
  wire[15:0] T234;
  wire[15:0] T235;
  wire[15:0] T236;
  wire[11:0] T237;
  wire[15:0] T238;
  wire[15:0] T239;
  wire[15:0] T240;
  wire[7:0] T241;
  wire[15:0] T242;
  wire[15:0] T243;
  wire[15:0] T550;
  wire[7:0] T244;
  wire[15:0] T245;
  wire[15:0] T551;
  wire[11:0] T246;
  wire[15:0] T247;
  wire[15:0] T552;
  wire[13:0] T248;
  wire[15:0] T249;
  wire[15:0] T553;
  wire[14:0] T250;
  wire[26:0] T251;
  wire[26:0] T554;
  wire T252;
  wire[27:0] sigX3;
  wire[42:0] T253;
  wire T254;
  wire T255;
  wire[15:0] T256;
  wire[15:0] absSigSumExtraMask;
  wire[14:0] T257;
  wire[6:0] T258;
  wire[2:0] T259;
  wire T260;
  wire[2:0] T261;
  wire[6:0] T262;
  wire[14:0] T263;
  wire[16:0] T264;
  wire[3:0] normTo2ShiftDist;
  wire[3:0] estNormDist_5;
  wire[3:0] T265;
  wire[1:0] T266;
  wire T267;
  wire[1:0] T268;
  wire T269;
  wire[3:0] T270;
  wire[1:0] T271;
  wire T272;
  wire[1:0] T273;
  wire[3:0] T274;
  wire T275;
  wire[1:0] T276;
  wire T277;
  wire[1:0] T278;
  wire T279;
  wire[7:0] T280;
  wire[7:0] T281;
  wire[7:0] T282;
  wire[6:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[7:0] T286;
  wire[5:0] T287;
  wire[7:0] T288;
  wire[7:0] T289;
  wire[7:0] T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T293;
  wire[7:0] T555;
  wire[3:0] T294;
  wire[7:0] T295;
  wire[7:0] T556;
  wire[5:0] T296;
  wire[7:0] T297;
  wire[7:0] T557;
  wire[6:0] T298;
  wire[15:0] T299;
  wire[42:0] cFirstNormAbsSigSum;
  wire[42:0] T558;
  wire[41:0] T300;
  wire[41:0] notCDom_pos_firstNormAbsSigSum;
  wire[41:0] T301;
  wire[41:0] T302;
  wire[31:0] T303;
  wire[31:0] T559;
  wire[9:0] T304;
  wire[41:0] T560;
  wire[33:0] T305;
  wire T306;
  wire T307;
  wire[1:0] firstReduceSigSum;
  wire T308;
  wire[17:0] T309;
  wire T310;
  wire[15:0] T311;
  wire T312;
  wire T313;
  wire[1:0] firstReduceNotSigSum;
  wire T314;
  wire[17:0] T315;
  wire[74:0] notSigSum;
  wire T316;
  wire[15:0] T317;
  wire[32:0] T318;
  wire T319;
  wire[41:0] T320;
  wire[41:0] T321;
  wire[41:0] T322;
  wire[15:0] T323;
  wire[15:0] T561;
  wire[25:0] T324;
  wire T325;
  wire T326;
  wire[41:0] CDom_firstNormAbsSigSum;
  wire[41:0] T327;
  wire[41:0] T328;
  wire[41:0] T329;
  wire T330;
  wire[40:0] T331;
  wire[41:0] T562;
  wire T332;
  wire T333;
  wire T334;
  wire[41:0] T335;
  wire[41:0] T336;
  wire[41:0] T337;
  wire T338;
  wire[40:0] T339;
  wire[41:0] T563;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[41:0] T344;
  wire[41:0] T345;
  wire[41:0] T346;
  wire T347;
  wire[40:0] T348;
  wire[41:0] T564;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire[41:0] T353;
  wire[41:0] T354;
  wire T355;
  wire[40:0] T356;
  wire[41:0] T565;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire[42:0] T362;
  wire[42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[42:0] T363;
  wire[42:0] T364;
  wire[10:0] T365;
  wire[42:0] T566;
  wire[32:0] T366;
  wire T367;
  wire[31:0] T368;
  wire T369;
  wire[42:0] T370;
  wire[42:0] T567;
  wire[41:0] T371;
  wire[42:0] T372;
  wire[26:0] T373;
  wire T374;
  wire T375;
  wire[42:0] T568;
  wire T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[41:0] T380;
  wire[41:0] T381;
  wire roundPosBit;
  wire[27:0] T382;
  wire[27:0] T569;
  wire[26:0] roundPosMask;
  wire[26:0] T570;
  wire[25:0] T383;
  wire[25:0] T384;
  wire T385;
  wire allRound;
  wire allRoundExtra;
  wire[27:0] T386;
  wire[27:0] T571;
  wire[25:0] T387;
  wire[27:0] T388;
  wire doIncrSig;
  wire T389;
  wire T390;
  wire T391;
  wire commonCase;
  wire T392;
  wire notSpecial_addZeros;
  wire T393;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T394;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T395;
  wire isSpecialA;
  wire[1:0] T396;
  wire underflow;
  wire underflowY;
  wire T397;
  wire T398;
  wire[9:0] T572;
  wire[7:0] T399;
  wire sigX3Shift1;
  wire[1:0] T400;
  wire T401;
  wire overflow;
  wire overflowY;
  wire[2:0] T402;
  wire[10:0] sExpY;
  wire[10:0] T403;
  wire[10:0] T404;
  wire T405;
  wire[1:0] T406;
  wire[25:0] sigY3;
  wire[25:0] T407;
  wire[25:0] T408;
  wire[25:0] T409;
  wire[25:0] T410;
  wire[25:0] roundUp_sigY3;
  wire[25:0] T411;
  wire[25:0] T412;
  wire[27:0] T413;
  wire[27:0] T573;
  wire roundEven;
  wire T414;
  wire T415;
  wire T416;
  wire roundingMode_nearest_even;
  wire T417;
  wire T418;
  wire T419;
  wire[25:0] T420;
  wire[25:0] T421;
  wire roundUp;
  wire T422;
  wire T423;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T424;
  wire doNegSignSum;
  wire T425;
  wire T426;
  wire T427;
  wire isZeroY;
  wire[2:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire[25:0] T442;
  wire[25:0] T443;
  wire[27:0] T444;
  wire[27:0] T574;
  wire[26:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[10:0] T449;
  wire[10:0] T450;
  wire T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire[1:0] T455;
  wire invalid;
  wire notSigNaN_invalid;
  wire T456;
  wire T457;
  wire isInfC;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire isInfB;
  wire T462;
  wire T463;
  wire isInfA;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire isNaNB;
  wire T468;
  wire T469;
  wire isNaNA;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire isSigNaNC;
  wire T475;
  wire T476;
  wire isNaNC;
  wire T477;
  wire T478;
  wire isSigNaNB;
  wire T479;
  wire T480;
  wire isSigNaNA;
  wire T481;
  wire T482;
  wire[32:0] T483;
  wire[31:0] T484;
  wire[22:0] fractOut;
  wire[22:0] T485;
  wire[22:0] T575;
  wire T486;
  wire isSatOut;
  wire T487;
  wire overflowY_roundMagUp;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire isNaNOut;
  wire T492;
  wire T493;
  wire[22:0] fractY;
  wire[22:0] T494;
  wire[22:0] T495;
  wire[8:0] expOut;
  wire[8:0] T496;
  wire[8:0] T497;
  wire[8:0] T498;
  wire notNaN_isInfOut;
  wire T499;
  wire T500;
  wire T501;
  wire[8:0] T502;
  wire[8:0] T503;
  wire[8:0] T504;
  wire[8:0] T505;
  wire[8:0] T506;
  wire[8:0] T507;
  wire[8:0] T508;
  wire[8:0] T509;
  wire[8:0] T510;
  wire[8:0] T511;
  wire[8:0] T512;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T513;
  wire[8:0] T514;
  wire T515;
  wire T516;
  wire[8:0] expY;
  wire signOut;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;


  assign io_exceptionFlags = T0;
  assign T0 = {T455, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T385 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 28'h0;
  assign T4 = sigX3 & T529;
  assign T529 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T251 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T530;
  assign T530 = {24'h0, T8};
  assign T8 = sigX3[5'h1a:5'h1a];
  assign T9 = {T226, T10};
  assign T10 = {T207, T11};
  assign T11 = T12[4'h8:4'h8];
  assign T12 = T13[5'h18:5'h10];
  assign T13 = T14[8'h83:7'h6b];
  assign T14 = $signed(1025'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T15;
  assign T15 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'h9:1'h0];
  assign sExpX3 = sExpSum - T531;
  assign T531 = {4'h0, estNormDist};
  assign estNormDist = isCDominant ? CDom_estNormDist : T16;
  assign T16 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = T197 ? 7'h18 : T17;
  assign T17 = T196 ? 7'h19 : T18;
  assign T18 = T195 ? 7'h1a : T19;
  assign T19 = T194 ? 7'h1b : T20;
  assign T20 = T193 ? 7'h1c : T21;
  assign T21 = T192 ? 7'h1d : T22;
  assign T22 = T191 ? 7'h1e : T23;
  assign T23 = T190 ? 7'h1f : T24;
  assign T24 = T189 ? 7'h20 : T25;
  assign T25 = T188 ? 7'h21 : T26;
  assign T26 = T187 ? 7'h22 : T27;
  assign T27 = T186 ? 7'h23 : T28;
  assign T28 = T185 ? 7'h24 : T29;
  assign T29 = T184 ? 7'h25 : T30;
  assign T30 = T183 ? 7'h26 : T31;
  assign T31 = T182 ? 7'h27 : T32;
  assign T32 = T181 ? 7'h28 : T33;
  assign T33 = T180 ? 7'h29 : T34;
  assign T34 = T179 ? 7'h2a : T35;
  assign T35 = T178 ? 7'h2b : T36;
  assign T36 = T177 ? 7'h2c : T37;
  assign T37 = T176 ? 7'h2d : T38;
  assign T38 = T175 ? 7'h2e : T39;
  assign T39 = T174 ? 7'h2f : T40;
  assign T40 = T173 ? 7'h30 : T41;
  assign T41 = T172 ? 7'h31 : T42;
  assign T42 = T171 ? 7'h32 : T43;
  assign T43 = T170 ? 7'h33 : T44;
  assign T44 = T169 ? 7'h34 : T45;
  assign T45 = T168 ? 7'h35 : T46;
  assign T46 = T167 ? 7'h36 : T47;
  assign T47 = T166 ? 7'h37 : T48;
  assign T48 = T165 ? 7'h38 : T49;
  assign T49 = T164 ? 7'h39 : T50;
  assign T50 = T163 ? 7'h3a : T51;
  assign T51 = T162 ? 7'h3b : T52;
  assign T52 = T161 ? 7'h3c : T53;
  assign T53 = T160 ? 7'h3d : T54;
  assign T54 = T159 ? 7'h3e : T55;
  assign T55 = T158 ? 7'h3f : T56;
  assign T56 = T157 ? 7'h40 : T57;
  assign T57 = T156 ? 7'h41 : T58;
  assign T58 = T155 ? 7'h42 : T59;
  assign T59 = T154 ? 7'h43 : T60;
  assign T60 = T153 ? 7'h44 : T61;
  assign T61 = T152 ? 7'h45 : T62;
  assign T62 = T151 ? 7'h46 : T63;
  assign T63 = T150 ? 7'h47 : T64;
  assign T64 = T65 ? 7'h48 : 7'h49;
  assign T65 = T66[1'h1:1'h1];
  assign T66 = T544 ^ T67;
  assign T67 = T68 << 1'h1;
  assign T68 = 50'h0 | T69;
  assign T69 = sigSum[6'h32:1'h1];
  assign sigSum = T543 + alignedNegSigC;
  assign alignedNegSigC = T70[7'h4a:1'h0];
  assign T70 = {T139, T71};
  assign T71 = T76 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T73 ^ T72;
  assign T72 = io_op[1'h0:1'h0];
  assign T73 = io_c[6'h20:6'h20];
  assign signProd = T75 ^ T74;
  assign T74 = io_op[1'h1:1'h1];
  assign T75 = signA ^ signB;
  assign signB = io_b[6'h20:6'h20];
  assign signA = io_a[6'h20:6'h20];
  assign T76 = T77 != 24'h0;
  assign T77 = sigC & CExtraMask;
  assign CExtraMask = {T112, T78};
  assign T78 = T110 | T79;
  assign T79 = T80 & 8'haa;
  assign T80 = T81 << 1'h1;
  assign T81 = T82[3'h6:1'h0];
  assign T82 = T108 | T83;
  assign T83 = T84 & 8'hcc;
  assign T84 = T85 << 2'h2;
  assign T85 = T86[3'h5:1'h0];
  assign T86 = T106 | T87;
  assign T87 = T88 & 8'hf0;
  assign T88 = T89 << 3'h4;
  assign T89 = T90[2'h3:1'h0];
  assign T90 = T91[5'h17:5'h10];
  assign T91 = T92[7'h4d:6'h36];
  assign T92 = $signed(129'h100000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = T93[3'h6:1'h0];
  assign T93 = CAlignDist_floor ? 11'h0 : T94;
  assign T94 = T101 ? sNatCAlignDist : 11'h4a;
  assign sNatCAlignDist = sExpAlignedProd - T532;
  assign T532 = {2'h0, expC};
  assign expC = io_c[5'h1f:5'h17];
  assign sExpAlignedProd = T95 + 11'h1b;
  assign T95 = T96 + T533;
  assign T533 = {2'h0, expA};
  assign expA = io_a[5'h1f:5'h17];
  assign T96 = {T98, T97};
  assign T97 = expB[3'h7:1'h0];
  assign expB = io_b[5'h1f:5'h17];
  assign T98 = 3'h0 - T534;
  assign T534 = {2'h0, T99};
  assign T99 = T100 ^ 1'h1;
  assign T100 = expB[4'h8:4'h8];
  assign T101 = T102 < 10'h4a;
  assign T102 = sNatCAlignDist[4'h9:1'h0];
  assign CAlignDist_floor = isZeroProd | T103;
  assign T103 = sNatCAlignDist[4'ha:4'ha];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T104 == 3'h0;
  assign T104 = expB[4'h8:3'h6];
  assign isZeroA = T105 == 3'h0;
  assign T105 = expA[4'h8:3'h6];
  assign T106 = T535 & 8'hf;
  assign T535 = {4'h0, T107};
  assign T107 = T90 >> 3'h4;
  assign T108 = T536 & 8'h33;
  assign T536 = {2'h0, T109};
  assign T109 = T86 >> 2'h2;
  assign T110 = T537 & 8'h55;
  assign T537 = {1'h0, T111};
  assign T111 = T82 >> 1'h1;
  assign T112 = T135 | T113;
  assign T113 = T114 & 16'haaaa;
  assign T114 = T115 << 1'h1;
  assign T115 = T116[4'he:1'h0];
  assign T116 = T133 | T117;
  assign T117 = T118 & 16'hcccc;
  assign T118 = T119 << 2'h2;
  assign T119 = T120[4'hd:1'h0];
  assign T120 = T131 | T121;
  assign T121 = T122 & 16'hf0f0;
  assign T122 = T123 << 3'h4;
  assign T123 = T124[4'hb:1'h0];
  assign T124 = T129 | T125;
  assign T125 = T126 & 16'hff00;
  assign T126 = T127 << 4'h8;
  assign T127 = T128[3'h7:1'h0];
  assign T128 = T91[4'hf:1'h0];
  assign T129 = T538 & 16'hff;
  assign T538 = {8'h0, T130};
  assign T130 = T128 >> 4'h8;
  assign T131 = T539 & 16'hf0f;
  assign T539 = {4'h0, T132};
  assign T132 = T124 >> 3'h4;
  assign T133 = T540 & 16'h3333;
  assign T540 = {2'h0, T134};
  assign T134 = T120 >> 2'h2;
  assign T135 = T541 & 16'h5555;
  assign T541 = {1'h0, T136};
  assign T136 = T116 >> 1'h1;
  assign sigC = {T137, fractC};
  assign fractC = io_c[5'h16:1'h0];
  assign T137 = isZeroC ^ 1'h1;
  assign isZeroC = T138 == 3'h0;
  assign T138 = expC[4'h8:3'h6];
  assign T139 = $signed(T140) >>> CAlignDist;
  assign T140 = T141;
  assign T141 = {doSubMags, T142};
  assign T142 = {negSigC, T143};
  assign T143 = 50'h0 - T542;
  assign T542 = {49'h0, doSubMags};
  assign negSigC = doSubMags ? T144 : sigC;
  assign T144 = ~ sigC;
  assign T543 = {26'h0, T145};
  assign T145 = T146 << 1'h1;
  assign T146 = sigA * sigB;
  assign sigB = {T147, fractB};
  assign fractB = io_b[5'h16:1'h0];
  assign T147 = isZeroB ^ 1'h1;
  assign sigA = {T148, fractA};
  assign fractA = io_a[5'h16:1'h0];
  assign T148 = isZeroA ^ 1'h1;
  assign T544 = {1'h0, T149};
  assign T149 = 50'h0 ^ T69;
  assign T150 = T66[2'h2:2'h2];
  assign T151 = T66[2'h3:2'h3];
  assign T152 = T66[3'h4:3'h4];
  assign T153 = T66[3'h5:3'h5];
  assign T154 = T66[3'h6:3'h6];
  assign T155 = T66[3'h7:3'h7];
  assign T156 = T66[4'h8:4'h8];
  assign T157 = T66[4'h9:4'h9];
  assign T158 = T66[4'ha:4'ha];
  assign T159 = T66[4'hb:4'hb];
  assign T160 = T66[4'hc:4'hc];
  assign T161 = T66[4'hd:4'hd];
  assign T162 = T66[4'he:4'he];
  assign T163 = T66[4'hf:4'hf];
  assign T164 = T66[5'h10:5'h10];
  assign T165 = T66[5'h11:5'h11];
  assign T166 = T66[5'h12:5'h12];
  assign T167 = T66[5'h13:5'h13];
  assign T168 = T66[5'h14:5'h14];
  assign T169 = T66[5'h15:5'h15];
  assign T170 = T66[5'h16:5'h16];
  assign T171 = T66[5'h17:5'h17];
  assign T172 = T66[5'h18:5'h18];
  assign T173 = T66[5'h19:5'h19];
  assign T174 = T66[5'h1a:5'h1a];
  assign T175 = T66[5'h1b:5'h1b];
  assign T176 = T66[5'h1c:5'h1c];
  assign T177 = T66[5'h1d:5'h1d];
  assign T178 = T66[5'h1e:5'h1e];
  assign T179 = T66[5'h1f:5'h1f];
  assign T180 = T66[6'h20:6'h20];
  assign T181 = T66[6'h21:6'h21];
  assign T182 = T66[6'h22:6'h22];
  assign T183 = T66[6'h23:6'h23];
  assign T184 = T66[6'h24:6'h24];
  assign T185 = T66[6'h25:6'h25];
  assign T186 = T66[6'h26:6'h26];
  assign T187 = T66[6'h27:6'h27];
  assign T188 = T66[6'h28:6'h28];
  assign T189 = T66[6'h29:6'h29];
  assign T190 = T66[6'h2a:6'h2a];
  assign T191 = T66[6'h2b:6'h2b];
  assign T192 = T66[6'h2c:6'h2c];
  assign T193 = T66[6'h2d:6'h2d];
  assign T194 = T66[6'h2e:6'h2e];
  assign T195 = T66[6'h2f:6'h2f];
  assign T196 = T66[6'h30:6'h30];
  assign T197 = T66[6'h31:6'h31];
  assign notCDom_signSigSum = sigSum[6'h33:6'h33];
  assign CDom_estNormDist = T200 ? CAlignDist : T545;
  assign T545 = {2'h0, T198};
  assign T198 = T199[3'h4:1'h0];
  assign T199 = CAlignDist - 7'h1;
  assign T200 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T201;
  assign T201 = T202 == 10'h0;
  assign T202 = sNatCAlignDist[4'h9:1'h0];
  assign isCDominant = T206 & T203;
  assign T203 = CAlignDist_floor | T204;
  assign T204 = T205 < 10'h19;
  assign T205 = sNatCAlignDist[4'h9:1'h0];
  assign T206 = isZeroC ^ 1'h1;
  assign sExpSum = CAlignDist_floor ? T546 : sExpAlignedProd;
  assign T546 = {2'h0, expC};
  assign T207 = T224 | T208;
  assign T208 = T209 & 8'haa;
  assign T209 = T210 << 1'h1;
  assign T210 = T211[3'h6:1'h0];
  assign T211 = T222 | T212;
  assign T212 = T213 & 8'hcc;
  assign T213 = T214 << 2'h2;
  assign T214 = T215[3'h5:1'h0];
  assign T215 = T220 | T216;
  assign T216 = T217 & 8'hf0;
  assign T217 = T218 << 3'h4;
  assign T218 = T219[2'h3:1'h0];
  assign T219 = T12[3'h7:1'h0];
  assign T220 = T547 & 8'hf;
  assign T547 = {4'h0, T221};
  assign T221 = T219 >> 3'h4;
  assign T222 = T548 & 8'h33;
  assign T548 = {2'h0, T223};
  assign T223 = T215 >> 2'h2;
  assign T224 = T549 & 8'h55;
  assign T549 = {1'h0, T225};
  assign T225 = T211 >> 1'h1;
  assign T226 = T249 | T227;
  assign T227 = T228 & 16'haaaa;
  assign T228 = T229 << 1'h1;
  assign T229 = T230[4'he:1'h0];
  assign T230 = T247 | T231;
  assign T231 = T232 & 16'hcccc;
  assign T232 = T233 << 2'h2;
  assign T233 = T234[4'hd:1'h0];
  assign T234 = T245 | T235;
  assign T235 = T236 & 16'hf0f0;
  assign T236 = T237 << 3'h4;
  assign T237 = T238[4'hb:1'h0];
  assign T238 = T243 | T239;
  assign T239 = T240 & 16'hff00;
  assign T240 = T241 << 4'h8;
  assign T241 = T242[3'h7:1'h0];
  assign T242 = T13[4'hf:1'h0];
  assign T243 = T550 & 16'hff;
  assign T550 = {8'h0, T244};
  assign T244 = T242 >> 4'h8;
  assign T245 = T551 & 16'hf0f;
  assign T551 = {4'h0, T246};
  assign T246 = T238 >> 3'h4;
  assign T247 = T552 & 16'h3333;
  assign T552 = {2'h0, T248};
  assign T248 = T234 >> 2'h2;
  assign T249 = T553 & 16'h5555;
  assign T553 = {1'h0, T250};
  assign T250 = T230 >> 1'h1;
  assign T251 = 27'h0 - T554;
  assign T554 = {26'h0, T252};
  assign T252 = sExpX3[4'ha:4'ha];
  assign sigX3 = T253[5'h1b:1'h0];
  assign T253 = {T380, T254};
  assign T254 = doIncrSig ? T376 : T255;
  assign T255 = T256 != 16'h0;
  assign T256 = T299 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T257, 1'h1};
  assign T257 = {T280, T258};
  assign T258 = {T270, T259};
  assign T259 = {T266, T260};
  assign T260 = T261[2'h2:2'h2];
  assign T261 = T262[3'h6:3'h4];
  assign T262 = T263[4'he:4'h8];
  assign T263 = T264[4'hf:1'h1];
  assign T264 = $signed(17'h10000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T265;
  assign T265 = estNormDist[2'h3:1'h0];
  assign T266 = {T269, T267};
  assign T267 = T268[1'h1:1'h1];
  assign T268 = T261[1'h1:1'h0];
  assign T269 = T268[1'h0:1'h0];
  assign T270 = {T276, T271};
  assign T271 = {T275, T272};
  assign T272 = T273[1'h1:1'h1];
  assign T273 = T274[2'h3:2'h2];
  assign T274 = T262[2'h3:1'h0];
  assign T275 = T273[1'h0:1'h0];
  assign T276 = {T279, T277};
  assign T277 = T278[1'h1:1'h1];
  assign T278 = T274[1'h1:1'h0];
  assign T279 = T278[1'h0:1'h0];
  assign T280 = T297 | T281;
  assign T281 = T282 & 8'haa;
  assign T282 = T283 << 1'h1;
  assign T283 = T284[3'h6:1'h0];
  assign T284 = T295 | T285;
  assign T285 = T286 & 8'hcc;
  assign T286 = T287 << 2'h2;
  assign T287 = T288[3'h5:1'h0];
  assign T288 = T293 | T289;
  assign T289 = T290 & 8'hf0;
  assign T290 = T291 << 3'h4;
  assign T291 = T292[2'h3:1'h0];
  assign T292 = T263[3'h7:1'h0];
  assign T293 = T555 & 8'hf;
  assign T555 = {4'h0, T294};
  assign T294 = T292 >> 3'h4;
  assign T295 = T556 & 8'h33;
  assign T556 = {2'h0, T296};
  assign T296 = T288 >> 2'h2;
  assign T297 = T557 & 8'h55;
  assign T557 = {1'h0, T298};
  assign T298 = T284 >> 1'h1;
  assign T299 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T362 : T558;
  assign T558 = {1'h0, T300};
  assign T300 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T326 ? T320 : T301;
  assign T301 = T319 ? T560 : T302;
  assign T302 = {T304, T303};
  assign T303 = 32'h0 - T559;
  assign T559 = {31'h0, doSubMags};
  assign T304 = sigSum[4'ha:1'h1];
  assign T560 = {8'h0, T305};
  assign T305 = {T318, T306};
  assign T306 = doSubMags ? T312 : T307;
  assign T307 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T310, T308};
  assign T308 = T309 != 18'h0;
  assign T309 = sigSum[5'h11:1'h0];
  assign T310 = T311 != 16'h0;
  assign T311 = sigSum[6'h21:5'h12];
  assign T312 = ~ T313;
  assign T313 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T316, T314};
  assign T314 = T315 != 18'h0;
  assign T315 = notSigSum[5'h11:1'h0];
  assign notSigSum = ~ sigSum;
  assign T316 = T317 != 16'h0;
  assign T317 = notSigSum[6'h21:5'h12];
  assign T318 = sigSum[6'h32:5'h12];
  assign T319 = estNormNeg_dist[3'h4:3'h4];
  assign T320 = T325 ? T322 : T321;
  assign T321 = sigSum[6'h2a:1'h1];
  assign T322 = {T324, T323};
  assign T323 = 16'h0 - T561;
  assign T561 = {15'h0, doSubMags};
  assign T324 = sigSum[5'h1a:1'h1];
  assign T325 = estNormNeg_dist[3'h4:3'h4];
  assign T326 = estNormNeg_dist[3'h5:3'h5];
  assign CDom_firstNormAbsSigSum = T327;
  assign T327 = T335 | T328;
  assign T328 = T562 & T329;
  assign T329 = {T331, T330};
  assign T330 = firstReduceNotSigSum[1'h0:1'h0];
  assign T331 = notSigSum[6'h3a:5'h12];
  assign T562 = T332 ? 42'h3ffffffffff : 42'h0;
  assign T332 = T333;
  assign T333 = doSubMags & T334;
  assign T334 = CDom_estNormDist[3'h4:3'h4];
  assign T335 = T344 | T336;
  assign T336 = T563 & T337;
  assign T337 = {T339, T338};
  assign T338 = firstReduceNotSigSum != 2'h0;
  assign T339 = notSigSum[7'h4a:6'h22];
  assign T563 = T340 ? 42'h3ffffffffff : 42'h0;
  assign T340 = T341;
  assign T341 = doSubMags & T342;
  assign T342 = ~ T343;
  assign T343 = CDom_estNormDist[3'h4:3'h4];
  assign T344 = T353 | T345;
  assign T345 = T564 & T346;
  assign T346 = {T348, T347};
  assign T347 = firstReduceSigSum[1'h0:1'h0];
  assign T348 = sigSum[6'h3a:5'h12];
  assign T564 = T349 ? 42'h3ffffffffff : 42'h0;
  assign T349 = T350;
  assign T350 = T352 & T351;
  assign T351 = CDom_estNormDist[3'h4:3'h4];
  assign T352 = ~ doSubMags;
  assign T353 = T565 & T354;
  assign T354 = {T356, T355};
  assign T355 = firstReduceSigSum != 2'h0;
  assign T356 = sigSum[7'h4a:6'h22];
  assign T565 = T357 ? 42'h3ffffffffff : 42'h0;
  assign T357 = T358;
  assign T358 = T361 & T359;
  assign T359 = ~ T360;
  assign T360 = CDom_estNormDist[3'h4:3'h4];
  assign T361 = ~ doSubMags;
  assign T362 = isCDominant ? T568 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T375 ? T370 : T363;
  assign T363 = T369 ? T566 : T364;
  assign T364 = T365 << 6'h20;
  assign T365 = notSigSum[4'hb:1'h1];
  assign T566 = {10'h0, T366};
  assign T366 = {T368, T367};
  assign T367 = firstReduceNotSigSum[1'h0:1'h0];
  assign T368 = notSigSum[6'h31:5'h12];
  assign T369 = estNormNeg_dist[3'h4:3'h4];
  assign T370 = T374 ? T372 : T567;
  assign T567 = {1'h0, T371};
  assign T371 = notSigSum[6'h2a:1'h1];
  assign T372 = T373 << 5'h10;
  assign T373 = notSigSum[5'h1b:1'h1];
  assign T374 = estNormNeg_dist[3'h4:3'h4];
  assign T375 = estNormNeg_dist[3'h5:3'h5];
  assign T568 = {1'h0, CDom_firstNormAbsSigSum};
  assign T376 = T377 == 16'h0;
  assign T377 = T378 & absSigSumExtraMask;
  assign T378 = ~ T379;
  assign T379 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign T380 = T381 >> normTo2ShiftDist;
  assign T381 = cFirstNormAbsSigSum[6'h2a:1'h1];
  assign roundPosBit = T382 != 28'h0;
  assign T382 = sigX3 & T569;
  assign T569 = {1'h0, roundPosMask};
  assign roundPosMask = T570 & roundMask;
  assign T570 = {1'h0, T383};
  assign T383 = ~ T384;
  assign T384 = roundMask >> 1'h1;
  assign T385 = ~ allRound;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T386 == 28'h0;
  assign T386 = T388 & T571;
  assign T571 = {2'h0, T387};
  assign T387 = roundMask >> 1'h1;
  assign T388 = ~ sigX3;
  assign doIncrSig = T389 & doSubMags;
  assign T389 = T391 & T390;
  assign T390 = ~ notCDom_signSigSum;
  assign T391 = ~ isCDominant;
  assign commonCase = T393 & T392;
  assign T392 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T393 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T394 == 2'h3;
  assign T394 = expC[4'h8:3'h7];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T395 == 2'h3;
  assign T395 = expB[4'h8:3'h7];
  assign isSpecialA = T396 == 2'h3;
  assign T396 = expA[4'h8:3'h7];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T397;
  assign T397 = T401 | T398;
  assign T398 = sExpX3_13 <= T572;
  assign T572 = {2'h0, T399};
  assign T399 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign sigX3Shift1 = T400 == 2'h0;
  assign T400 = sigX3[5'h1b:5'h1a];
  assign T401 = sExpX3[4'ha:4'ha];
  assign overflow = commonCase & overflowY;
  assign overflowY = T402 == 3'h3;
  assign T402 = sExpY[4'h9:3'h7];
  assign sExpY = T449 | T403;
  assign T403 = T405 ? T404 : 11'h0;
  assign T404 = sExpX3 - 11'h1;
  assign T405 = T406 == 2'h0;
  assign T406 = sigY3[5'h19:5'h18];
  assign sigY3 = T420 | T407;
  assign T407 = roundEven ? T408 : 26'h0;
  assign T408 = roundUp_sigY3 & T409;
  assign T409 = ~ T410;
  assign T410 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T411[5'h19:1'h0];
  assign T411 = T412 + 26'h1;
  assign T412 = T413 >> 2'h2;
  assign T413 = sigX3 | T573;
  assign T573 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T417 : T414;
  assign T414 = T416 & T415;
  assign T415 = ~ anyRoundExtra;
  assign T416 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T417 = T418 & allRoundExtra;
  assign T418 = roundingMode_nearest_even & T419;
  assign T419 = ~ roundPosBit;
  assign T420 = T442 | T421;
  assign T421 = roundUp ? roundUp_sigY3 : 26'h0;
  assign roundUp = T429 | T422;
  assign T422 = T423 & 1'h1;
  assign T423 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T427 & T424;
  assign T424 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T425 : notCDom_signSigSum;
  assign T425 = doSubMags & T426;
  assign T426 = ~ isZeroC;
  assign T427 = ~ isZeroY;
  assign isZeroY = T428 == 3'h0;
  assign T428 = sigX3[5'h1b:5'h19];
  assign T429 = T432 | T430;
  assign T430 = T431 & roundPosBit;
  assign T431 = doIncrSig & roundingMode_nearest_even;
  assign T432 = T434 | T433;
  assign T433 = doIncrSig & allRound;
  assign T434 = T438 | T435;
  assign T435 = T436 & anyRound;
  assign T436 = T437 & roundDirectUp;
  assign T437 = ~ doIncrSig;
  assign T438 = T439 & anyRoundExtra;
  assign T439 = T440 & roundPosBit;
  assign T440 = T441 & roundingMode_nearest_even;
  assign T441 = ~ doIncrSig;
  assign T442 = T446 ? T443 : 26'h0;
  assign T443 = T444 >> 2'h2;
  assign T444 = sigX3 & T574;
  assign T574 = {1'h0, T445};
  assign T445 = ~ roundMask;
  assign T446 = T448 & T447;
  assign T447 = ~ roundEven;
  assign T448 = ~ roundUp;
  assign T449 = T452 | T450;
  assign T450 = T451 ? sExpX3 : 11'h0;
  assign T451 = sigY3[5'h18:5'h18];
  assign T452 = T454 ? T453 : 11'h0;
  assign T453 = sExpX3 + 11'h1;
  assign T454 = sigY3[5'h19:5'h19];
  assign T455 = {invalid, 1'h0};
  assign invalid = T474 | notSigNaN_invalid;
  assign notSigNaN_invalid = T471 | T456;
  assign T456 = T457 & doSubMags;
  assign T457 = T460 & isInfC;
  assign isInfC = isSpecialC & T458;
  assign T458 = T459 ^ 1'h1;
  assign T459 = expC[3'h6:3'h6];
  assign T460 = T466 & T461;
  assign T461 = isInfA | isInfB;
  assign isInfB = isSpecialB & T462;
  assign T462 = T463 ^ 1'h1;
  assign T463 = expB[3'h6:3'h6];
  assign isInfA = isSpecialA & T464;
  assign T464 = T465 ^ 1'h1;
  assign T465 = expA[3'h6:3'h6];
  assign T466 = T469 & T467;
  assign T467 = ~ isNaNB;
  assign isNaNB = isSpecialB & T468;
  assign T468 = expB[3'h6:3'h6];
  assign T469 = ~ isNaNA;
  assign isNaNA = isSpecialA & T470;
  assign T470 = expA[3'h6:3'h6];
  assign T471 = T473 | T472;
  assign T472 = isZeroA & isInfB;
  assign T473 = isInfA & isZeroB;
  assign T474 = T478 | isSigNaNC;
  assign isSigNaNC = isNaNC & T475;
  assign T475 = T476 ^ 1'h1;
  assign T476 = fractC[5'h16:5'h16];
  assign isNaNC = isSpecialC & T477;
  assign T477 = expC[3'h6:3'h6];
  assign T478 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T479;
  assign T479 = T480 ^ 1'h1;
  assign T480 = fractB[5'h16:5'h16];
  assign isSigNaNA = isNaNA & T481;
  assign T481 = T482 ^ 1'h1;
  assign T482 = fractA[5'h16:5'h16];
  assign io_out = T483;
  assign T483 = {signOut, T484};
  assign T484 = {expOut, fractOut};
  assign fractOut = fractY | T485;
  assign T485 = 23'h0 - T575;
  assign T575 = {22'h0, T486};
  assign T486 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T487;
  assign T487 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T490 | T488;
  assign T488 = roundingMode_max & T489;
  assign T489 = ~ signY;
  assign T490 = roundingMode_nearest_even | T491;
  assign T491 = roundingMode_min & signY;
  assign isNaNOut = T492 | notSigNaN_invalid;
  assign T492 = T493 | isNaNC;
  assign T493 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T495 : T494;
  assign T494 = sigY3[5'h17:1'h1];
  assign T495 = sigY3[5'h16:1'h0];
  assign expOut = T497 | T496;
  assign T496 = isNaNOut ? 9'h1c0 : 9'h0;
  assign T497 = T502 | T498;
  assign T498 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign notNaN_isInfOut = T500 | T499;
  assign T499 = overflow & overflowY_roundMagUp;
  assign T500 = T501 | isInfC;
  assign T501 = isInfA | isInfB;
  assign T502 = T504 | T503;
  assign T503 = isSatOut ? 9'h17f : 9'h0;
  assign T504 = T507 & T505;
  assign T505 = ~ T506;
  assign T506 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T507 = T510 & T508;
  assign T508 = ~ T509;
  assign T509 = isSatOut ? 9'h80 : 9'h0;
  assign T510 = expY & T511;
  assign T511 = ~ T512;
  assign T512 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign notSpecial_isZeroOut = T516 | totalUnderflowY;
  assign totalUnderflowY = T515 | T513;
  assign T513 = T514 < 9'h6b;
  assign T514 = sExpY[4'h8:1'h0];
  assign T515 = sExpY[4'h9:4'h9];
  assign T516 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'h8:1'h0];
  assign signOut = T518 | T517;
  assign T517 = commonCase & signY;
  assign T518 = T522 | T519;
  assign T519 = T520 & opSignC;
  assign T520 = T521 & isSpecialC;
  assign T521 = mulSpecial ^ 1'h1;
  assign T522 = T526 | T523;
  assign T523 = T524 & signProd;
  assign T524 = mulSpecial & T525;
  assign T525 = isSpecialC ^ 1'h1;
  assign T526 = T527 | isNaNOut;
  assign T527 = T528 & opSignC;
  assign T528 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_0(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T25;
  reg [2:0] in_rm;
  wire[2:0] T0;
  wire[32:0] T26;
  reg [64:0] in_in3;
  wire[64:0] T1;
  wire[64:0] T2;
  wire[64:0] T27;
  wire[32:0] zero;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[32:0] T28;
  reg [64:0] in_in2;
  wire[64:0] T9;
  wire[64:0] T10;
  wire T11;
  wire[32:0] T29;
  reg [64:0] in_in1;
  wire[64:0] T12;
  wire[1:0] T30;
  reg [4:0] in_cmd;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[4:0] T31;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [4:0] R20;
  wire[4:0] T21;
  wire[4:0] res_exc;
  reg  valid;
  reg [64:0] R22;
  wire[64:0] T23;
  wire[64:0] res_data;
  wire[64:0] T32;
  reg  R24;
  wire T33;
  wire[32:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R20 = {1{$random}};
    valid = {1{$random}};
    R22 = {3{$random}};
    R24 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T25 = in_rm[1'h1:1'h0];
  assign T0 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T26 = in_in3[6'h20:1'h0];
  assign T1 = T6 ? T27 : T2;
  assign T2 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T27 = {32'h0, zero};
  assign zero = T3 << 6'h20;
  assign T3 = T5 ^ T4;
  assign T4 = io_in_bits_in2[6'h20:6'h20];
  assign T5 = io_in_bits_in1[6'h20:6'h20];
  assign T6 = io_in_valid & T7;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T28 = in_in2[6'h20:1'h0];
  assign T9 = T11 ? 65'h80000000 : T10;
  assign T10 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T11 = io_in_valid & io_in_bits_swap23;
  assign T29 = in_in1[6'h20:1'h0];
  assign T12 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T30 = in_cmd[1'h1:1'h0];
  assign T13 = io_in_valid ? T31 : T14;
  assign T14 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T31 = {3'h0, T15};
  assign T15 = {T17, T16};
  assign T16 = io_in_bits_cmd[1'h0:1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T19 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R20;
  assign T21 = valid ? res_exc : R20;
  assign res_exc = fma_io_exceptionFlags;
  assign io_out_bits_data = R22;
  assign T23 = valid ? res_data : R22;
  assign res_data = T32;
  assign T32 = {32'h0, fma_io_out};
  assign io_out_valid = R24;
  assign T33 = reset ? 1'h0 : valid;
  mulAddSubRecodedFloatN_0 fma(
       .io_op( T30 ),
       .io_a( T29 ),
       .io_b( T28 ),
       .io_c( T26 ),
       .io_roundingMode( T25 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T6) begin
      in_in3 <= T27;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T11) begin
      in_in2 <= 65'h80000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T31;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(valid) begin
      R20 <= res_exc;
    end
    valid <= io_in_valid;
    if(valid) begin
      R22 <= res_data;
    end
    if(reset) begin
      R24 <= 1'h0;
    end else begin
      R24 <= valid;
    end
  end
endmodule

module mulAddSubRecodedFloatN_1(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire inexactY;
  wire anyRound;
  wire anyRoundExtra;
  wire[56:0] T4;
  wire[56:0] T744;
  wire[54:0] T5;
  wire[55:0] roundMask;
  wire[55:0] T6;
  wire[53:0] T7;
  wire[53:0] T745;
  wire T8;
  wire[53:0] T9;
  wire[21:0] T10;
  wire[5:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[5:0] T15;
  wire[21:0] T16;
  wire[53:0] T17;
  wire[8192:0] T18;
  wire[12:0] T19;
  wire[12:0] sExpX3_13;
  wire[13:0] sExpX3;
  wire[13:0] T746;
  wire[7:0] estNormDist;
  wire[7:0] T20;
  wire[7:0] estNormNeg_dist;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire[7:0] T25;
  wire[7:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[7:0] T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[7:0] T58;
  wire[7:0] T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire[7:0] T75;
  wire[7:0] T76;
  wire[7:0] T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire[7:0] T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T119;
  wire[7:0] T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire T127;
  wire[108:0] T128;
  wire[108:0] T129;
  wire[107:0] T130;
  wire[107:0] T131;
  wire[161:0] sigSum;
  wire[161:0] alignedNegSigC;
  wire[162:0] T132;
  wire T133;
  wire doSubMags;
  wire opSignC;
  wire T134;
  wire T135;
  wire signProd;
  wire T136;
  wire T137;
  wire signB;
  wire signA;
  wire T138;
  wire[52:0] T139;
  wire[52:0] CExtraMask;
  wire[20:0] T140;
  wire[4:0] T141;
  wire T142;
  wire[4:0] T143;
  wire[20:0] T144;
  wire[52:0] T145;
  wire[256:0] T146;
  wire[7:0] CAlignDist;
  wire[13:0] T147;
  wire[13:0] T148;
  wire[13:0] sNatCAlignDist;
  wire[13:0] T747;
  wire[11:0] expC;
  wire[13:0] sExpAlignedProd;
  wire[13:0] T149;
  wire[13:0] T748;
  wire[11:0] expA;
  wire[13:0] T150;
  wire[10:0] T151;
  wire[11:0] expB;
  wire[2:0] T152;
  wire[2:0] T749;
  wire T153;
  wire T154;
  wire T155;
  wire[12:0] T156;
  wire CAlignDist_floor;
  wire T157;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T158;
  wire isZeroA;
  wire[2:0] T159;
  wire[3:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[1:0] T163;
  wire[3:0] T164;
  wire T165;
  wire[1:0] T166;
  wire T167;
  wire[1:0] T168;
  wire T169;
  wire[15:0] T170;
  wire[15:0] T171;
  wire[15:0] T172;
  wire[14:0] T173;
  wire[15:0] T174;
  wire[15:0] T175;
  wire[15:0] T176;
  wire[13:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[15:0] T180;
  wire[11:0] T181;
  wire[15:0] T182;
  wire[15:0] T183;
  wire[15:0] T184;
  wire[7:0] T185;
  wire[15:0] T186;
  wire[15:0] T187;
  wire[15:0] T750;
  wire[7:0] T188;
  wire[15:0] T189;
  wire[15:0] T751;
  wire[11:0] T190;
  wire[15:0] T191;
  wire[15:0] T752;
  wire[13:0] T192;
  wire[15:0] T193;
  wire[15:0] T753;
  wire[14:0] T194;
  wire[31:0] T195;
  wire[31:0] T196;
  wire[31:0] T197;
  wire[30:0] T198;
  wire[31:0] T199;
  wire[31:0] T200;
  wire[31:0] T201;
  wire[29:0] T202;
  wire[31:0] T203;
  wire[31:0] T204;
  wire[31:0] T205;
  wire[27:0] T206;
  wire[31:0] T207;
  wire[31:0] T208;
  wire[31:0] T209;
  wire[23:0] T210;
  wire[31:0] T211;
  wire[31:0] T212;
  wire[31:0] T213;
  wire[15:0] T214;
  wire[31:0] T215;
  wire[31:0] T216;
  wire[31:0] T754;
  wire[15:0] T217;
  wire[31:0] T218;
  wire[31:0] T755;
  wire[23:0] T219;
  wire[31:0] T220;
  wire[31:0] T756;
  wire[27:0] T221;
  wire[31:0] T222;
  wire[31:0] T757;
  wire[29:0] T223;
  wire[31:0] T224;
  wire[31:0] T758;
  wire[30:0] T225;
  wire[52:0] sigC;
  wire[51:0] fractC;
  wire T226;
  wire isZeroC;
  wire[2:0] T227;
  wire[161:0] T228;
  wire[161:0] T229;
  wire[161:0] T230;
  wire[160:0] T231;
  wire[107:0] T232;
  wire[107:0] T759;
  wire[52:0] negSigC;
  wire[52:0] T233;
  wire[161:0] T760;
  wire[106:0] T234;
  wire[105:0] T235;
  wire[52:0] sigB;
  wire[51:0] fractB;
  wire T236;
  wire[52:0] sigA;
  wire[51:0] fractA;
  wire T237;
  wire[108:0] T761;
  wire[107:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire notCDom_signSigSum;
  wire[7:0] CDom_estNormDist;
  wire[7:0] T762;
  wire[5:0] T345;
  wire[7:0] T346;
  wire T347;
  wire CAlignDist_0;
  wire T348;
  wire[12:0] T349;
  wire isCDominant;
  wire T350;
  wire T351;
  wire[12:0] T352;
  wire T353;
  wire[13:0] sExpSum;
  wire[13:0] T763;
  wire T354;
  wire[3:0] T355;
  wire[1:0] T356;
  wire T357;
  wire[1:0] T358;
  wire[3:0] T359;
  wire T360;
  wire[1:0] T361;
  wire T362;
  wire[1:0] T363;
  wire T364;
  wire[15:0] T365;
  wire[15:0] T366;
  wire[15:0] T367;
  wire[14:0] T368;
  wire[15:0] T369;
  wire[15:0] T370;
  wire[15:0] T371;
  wire[13:0] T372;
  wire[15:0] T373;
  wire[15:0] T374;
  wire[15:0] T375;
  wire[11:0] T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[7:0] T380;
  wire[15:0] T381;
  wire[15:0] T382;
  wire[15:0] T764;
  wire[7:0] T383;
  wire[15:0] T384;
  wire[15:0] T765;
  wire[11:0] T385;
  wire[15:0] T386;
  wire[15:0] T766;
  wire[13:0] T387;
  wire[15:0] T388;
  wire[15:0] T767;
  wire[14:0] T389;
  wire[31:0] T390;
  wire[31:0] T391;
  wire[31:0] T392;
  wire[30:0] T393;
  wire[31:0] T394;
  wire[31:0] T395;
  wire[31:0] T396;
  wire[29:0] T397;
  wire[31:0] T398;
  wire[31:0] T399;
  wire[31:0] T400;
  wire[27:0] T401;
  wire[31:0] T402;
  wire[31:0] T403;
  wire[31:0] T404;
  wire[23:0] T405;
  wire[31:0] T406;
  wire[31:0] T407;
  wire[31:0] T408;
  wire[15:0] T409;
  wire[31:0] T410;
  wire[31:0] T411;
  wire[31:0] T768;
  wire[15:0] T412;
  wire[31:0] T413;
  wire[31:0] T769;
  wire[23:0] T414;
  wire[31:0] T415;
  wire[31:0] T770;
  wire[27:0] T416;
  wire[31:0] T417;
  wire[31:0] T771;
  wire[29:0] T418;
  wire[31:0] T419;
  wire[31:0] T772;
  wire[30:0] T420;
  wire[55:0] T421;
  wire[55:0] T773;
  wire T422;
  wire[56:0] sigX3;
  wire[87:0] T423;
  wire T424;
  wire T425;
  wire[31:0] T426;
  wire[31:0] absSigSumExtraMask;
  wire[30:0] T427;
  wire[14:0] T428;
  wire[6:0] T429;
  wire[2:0] T430;
  wire T431;
  wire[2:0] T432;
  wire[6:0] T433;
  wire[14:0] T434;
  wire[30:0] T435;
  wire[32:0] T436;
  wire[4:0] normTo2ShiftDist;
  wire[4:0] estNormDist_5;
  wire[4:0] T437;
  wire[1:0] T438;
  wire T439;
  wire[1:0] T440;
  wire T441;
  wire[3:0] T442;
  wire[1:0] T443;
  wire T444;
  wire[1:0] T445;
  wire[3:0] T446;
  wire T447;
  wire[1:0] T448;
  wire T449;
  wire[1:0] T450;
  wire T451;
  wire[7:0] T452;
  wire[7:0] T453;
  wire[7:0] T454;
  wire[6:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[5:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[3:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T774;
  wire[3:0] T466;
  wire[7:0] T467;
  wire[7:0] T775;
  wire[5:0] T468;
  wire[7:0] T469;
  wire[7:0] T776;
  wire[6:0] T470;
  wire[15:0] T471;
  wire[15:0] T472;
  wire[15:0] T473;
  wire[14:0] T474;
  wire[15:0] T475;
  wire[15:0] T476;
  wire[15:0] T477;
  wire[13:0] T478;
  wire[15:0] T479;
  wire[15:0] T480;
  wire[15:0] T481;
  wire[11:0] T482;
  wire[15:0] T483;
  wire[15:0] T484;
  wire[15:0] T485;
  wire[7:0] T486;
  wire[15:0] T487;
  wire[15:0] T488;
  wire[15:0] T777;
  wire[7:0] T489;
  wire[15:0] T490;
  wire[15:0] T778;
  wire[11:0] T491;
  wire[15:0] T492;
  wire[15:0] T779;
  wire[13:0] T493;
  wire[15:0] T494;
  wire[15:0] T780;
  wire[14:0] T495;
  wire[31:0] T496;
  wire[87:0] cFirstNormAbsSigSum;
  wire[87:0] T781;
  wire[86:0] T497;
  wire[86:0] notCDom_pos_firstNormAbsSigSum;
  wire[86:0] T498;
  wire[86:0] T499;
  wire[53:0] T500;
  wire[53:0] T782;
  wire[32:0] T501;
  wire[86:0] T502;
  wire[86:0] T503;
  wire[85:0] T504;
  wire[85:0] T783;
  wire T505;
  wire[86:0] T784;
  wire[65:0] T506;
  wire T507;
  wire T508;
  wire[1:0] firstReduceSigSum;
  wire T509;
  wire[43:0] T510;
  wire T511;
  wire[31:0] T512;
  wire T513;
  wire T514;
  wire[1:0] firstReduceNotSigSum;
  wire T515;
  wire[43:0] T516;
  wire[161:0] notSigSum;
  wire T517;
  wire[31:0] T518;
  wire[64:0] T519;
  wire T520;
  wire T521;
  wire[86:0] T522;
  wire[86:0] T523;
  wire T524;
  wire T525;
  wire[10:0] T526;
  wire T527;
  wire[10:0] T528;
  wire[85:0] T529;
  wire[86:0] T530;
  wire[21:0] T531;
  wire[21:0] T785;
  wire[64:0] T532;
  wire T533;
  wire T534;
  wire[86:0] CDom_firstNormAbsSigSum;
  wire[86:0] T535;
  wire[86:0] T536;
  wire[86:0] T537;
  wire T538;
  wire[85:0] T539;
  wire[86:0] T786;
  wire T540;
  wire T541;
  wire T542;
  wire[86:0] T543;
  wire[86:0] T544;
  wire[86:0] T545;
  wire T546;
  wire[85:0] T547;
  wire[86:0] T787;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire[86:0] T552;
  wire[86:0] T553;
  wire[86:0] T554;
  wire T555;
  wire[85:0] T556;
  wire[86:0] T788;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire[86:0] T561;
  wire[86:0] T562;
  wire T563;
  wire[85:0] T564;
  wire[86:0] T789;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire[87:0] T570;
  wire[87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[87:0] T571;
  wire[87:0] T572;
  wire[33:0] T573;
  wire[87:0] T574;
  wire[87:0] T575;
  wire[1:0] T576;
  wire[87:0] T790;
  wire[64:0] T577;
  wire T578;
  wire[63:0] T579;
  wire T580;
  wire T581;
  wire[87:0] T582;
  wire[87:0] T583;
  wire T584;
  wire[10:0] T585;
  wire[86:0] T586;
  wire[87:0] T587;
  wire[65:0] T588;
  wire T589;
  wire T590;
  wire[87:0] T791;
  wire T591;
  wire[31:0] T592;
  wire[31:0] T593;
  wire[31:0] T594;
  wire[86:0] T595;
  wire[86:0] T596;
  wire roundPosBit;
  wire[56:0] T597;
  wire[56:0] T792;
  wire[55:0] roundPosMask;
  wire[55:0] T793;
  wire[54:0] T598;
  wire[54:0] T599;
  wire T600;
  wire allRound;
  wire allRoundExtra;
  wire[56:0] T601;
  wire[56:0] T794;
  wire[54:0] T602;
  wire[56:0] T603;
  wire doIncrSig;
  wire T604;
  wire T605;
  wire T606;
  wire commonCase;
  wire T607;
  wire notSpecial_addZeros;
  wire T608;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T609;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T610;
  wire isSpecialA;
  wire[1:0] T611;
  wire underflow;
  wire underflowY;
  wire T612;
  wire T613;
  wire[12:0] T795;
  wire[10:0] T614;
  wire sigX3Shift1;
  wire[1:0] T615;
  wire T616;
  wire overflow;
  wire overflowY;
  wire[2:0] T617;
  wire[13:0] sExpY;
  wire[13:0] T618;
  wire[13:0] T619;
  wire T620;
  wire[1:0] T621;
  wire[54:0] sigY3;
  wire[54:0] T622;
  wire[54:0] T623;
  wire[54:0] T624;
  wire[54:0] T625;
  wire[54:0] roundUp_sigY3;
  wire[54:0] T626;
  wire[54:0] T627;
  wire[56:0] T628;
  wire[56:0] T796;
  wire roundEven;
  wire T629;
  wire T630;
  wire T631;
  wire roundingMode_nearest_even;
  wire T632;
  wire T633;
  wire T634;
  wire[54:0] T635;
  wire[54:0] T636;
  wire roundUp;
  wire T637;
  wire T638;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T639;
  wire doNegSignSum;
  wire T640;
  wire T641;
  wire T642;
  wire isZeroY;
  wire[2:0] T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire[54:0] T657;
  wire[54:0] T658;
  wire[56:0] T659;
  wire[56:0] T797;
  wire[55:0] T660;
  wire T661;
  wire T662;
  wire T663;
  wire[13:0] T664;
  wire[13:0] T665;
  wire T666;
  wire[13:0] T667;
  wire[13:0] T668;
  wire T669;
  wire[1:0] T670;
  wire invalid;
  wire notSigNaN_invalid;
  wire T671;
  wire T672;
  wire isInfC;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire isInfB;
  wire T677;
  wire T678;
  wire isInfA;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire isNaNB;
  wire T683;
  wire T684;
  wire isNaNA;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire isSigNaNC;
  wire T690;
  wire T691;
  wire isNaNC;
  wire T692;
  wire T693;
  wire isSigNaNB;
  wire T694;
  wire T695;
  wire isSigNaNA;
  wire T696;
  wire T697;
  wire[64:0] T698;
  wire[63:0] T699;
  wire[51:0] fractOut;
  wire[51:0] T700;
  wire[51:0] T798;
  wire T701;
  wire isSatOut;
  wire T702;
  wire overflowY_roundMagUp;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire isNaNOut;
  wire T707;
  wire T708;
  wire[51:0] fractY;
  wire[51:0] T709;
  wire[51:0] T710;
  wire[11:0] expOut;
  wire[11:0] T711;
  wire[11:0] T712;
  wire[11:0] T713;
  wire notNaN_isInfOut;
  wire T714;
  wire T715;
  wire T716;
  wire[11:0] T717;
  wire[11:0] T718;
  wire[11:0] T719;
  wire[11:0] T720;
  wire[11:0] T721;
  wire[11:0] T722;
  wire[11:0] T723;
  wire[11:0] T724;
  wire[11:0] T725;
  wire[11:0] T726;
  wire[11:0] T727;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T728;
  wire[11:0] T729;
  wire T730;
  wire T731;
  wire[11:0] expY;
  wire signOut;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;


  assign io_exceptionFlags = T0;
  assign T0 = {T670, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & inexactY;
  assign inexactY = doIncrSig ? T600 : anyRound;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign anyRoundExtra = T4 != 57'h0;
  assign T4 = sigX3 & T744;
  assign T744 = {2'h0, T5};
  assign T5 = roundMask >> 1'h1;
  assign roundMask = T421 | T6;
  assign T6 = {T7, 2'h3};
  assign T7 = T9 | T745;
  assign T745 = {53'h0, T8};
  assign T8 = sigX3[6'h37:6'h37];
  assign T9 = {T390, T10};
  assign T10 = {T365, T11};
  assign T11 = {T355, T12};
  assign T12 = {T354, T13};
  assign T13 = T14[1'h1:1'h1];
  assign T14 = T15[3'h5:3'h4];
  assign T15 = T16[5'h15:5'h10];
  assign T16 = T17[6'h35:6'h20];
  assign T17 = T18[11'h403:10'h3ce];
  assign T18 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T19;
  assign T19 = ~ sExpX3_13;
  assign sExpX3_13 = sExpX3[4'hc:1'h0];
  assign sExpX3 = sExpSum - T746;
  assign T746 = {6'h0, estNormDist};
  assign estNormDist = isCDominant ? CDom_estNormDist : T20;
  assign T20 = notCDom_signSigSum ? estNormNeg_dist : estNormNeg_dist;
  assign estNormNeg_dist = T344 ? 8'h35 : T21;
  assign T21 = T343 ? 8'h36 : T22;
  assign T22 = T342 ? 8'h37 : T23;
  assign T23 = T341 ? 8'h38 : T24;
  assign T24 = T340 ? 8'h39 : T25;
  assign T25 = T339 ? 8'h3a : T26;
  assign T26 = T338 ? 8'h3b : T27;
  assign T27 = T337 ? 8'h3c : T28;
  assign T28 = T336 ? 8'h3d : T29;
  assign T29 = T335 ? 8'h3e : T30;
  assign T30 = T334 ? 8'h3f : T31;
  assign T31 = T333 ? 8'h40 : T32;
  assign T32 = T332 ? 8'h41 : T33;
  assign T33 = T331 ? 8'h42 : T34;
  assign T34 = T330 ? 8'h43 : T35;
  assign T35 = T329 ? 8'h44 : T36;
  assign T36 = T328 ? 8'h45 : T37;
  assign T37 = T327 ? 8'h46 : T38;
  assign T38 = T326 ? 8'h47 : T39;
  assign T39 = T325 ? 8'h48 : T40;
  assign T40 = T324 ? 8'h49 : T41;
  assign T41 = T323 ? 8'h4a : T42;
  assign T42 = T322 ? 8'h4b : T43;
  assign T43 = T321 ? 8'h4c : T44;
  assign T44 = T320 ? 8'h4d : T45;
  assign T45 = T319 ? 8'h4e : T46;
  assign T46 = T318 ? 8'h4f : T47;
  assign T47 = T317 ? 8'h50 : T48;
  assign T48 = T316 ? 8'h51 : T49;
  assign T49 = T315 ? 8'h52 : T50;
  assign T50 = T314 ? 8'h53 : T51;
  assign T51 = T313 ? 8'h54 : T52;
  assign T52 = T312 ? 8'h55 : T53;
  assign T53 = T311 ? 8'h56 : T54;
  assign T54 = T310 ? 8'h57 : T55;
  assign T55 = T309 ? 8'h58 : T56;
  assign T56 = T308 ? 8'h59 : T57;
  assign T57 = T307 ? 8'h5a : T58;
  assign T58 = T306 ? 8'h5b : T59;
  assign T59 = T305 ? 8'h5c : T60;
  assign T60 = T304 ? 8'h5d : T61;
  assign T61 = T303 ? 8'h5e : T62;
  assign T62 = T302 ? 8'h5f : T63;
  assign T63 = T301 ? 8'h60 : T64;
  assign T64 = T300 ? 8'h61 : T65;
  assign T65 = T299 ? 8'h62 : T66;
  assign T66 = T298 ? 8'h63 : T67;
  assign T67 = T297 ? 8'h64 : T68;
  assign T68 = T296 ? 8'h65 : T69;
  assign T69 = T295 ? 8'h66 : T70;
  assign T70 = T294 ? 8'h67 : T71;
  assign T71 = T293 ? 8'h68 : T72;
  assign T72 = T292 ? 8'h69 : T73;
  assign T73 = T291 ? 8'h6a : T74;
  assign T74 = T290 ? 8'h6b : T75;
  assign T75 = T289 ? 8'h6c : T76;
  assign T76 = T288 ? 8'h6d : T77;
  assign T77 = T287 ? 8'h6e : T78;
  assign T78 = T286 ? 8'h6f : T79;
  assign T79 = T285 ? 8'h70 : T80;
  assign T80 = T284 ? 8'h71 : T81;
  assign T81 = T283 ? 8'h72 : T82;
  assign T82 = T282 ? 8'h73 : T83;
  assign T83 = T281 ? 8'h74 : T84;
  assign T84 = T280 ? 8'h75 : T85;
  assign T85 = T279 ? 8'h76 : T86;
  assign T86 = T278 ? 8'h77 : T87;
  assign T87 = T277 ? 8'h78 : T88;
  assign T88 = T276 ? 8'h79 : T89;
  assign T89 = T275 ? 8'h7a : T90;
  assign T90 = T274 ? 8'h7b : T91;
  assign T91 = T273 ? 8'h7c : T92;
  assign T92 = T272 ? 8'h7d : T93;
  assign T93 = T271 ? 8'h7e : T94;
  assign T94 = T270 ? 8'h7f : T95;
  assign T95 = T269 ? 8'h80 : T96;
  assign T96 = T268 ? 8'h81 : T97;
  assign T97 = T267 ? 8'h82 : T98;
  assign T98 = T266 ? 8'h83 : T99;
  assign T99 = T265 ? 8'h84 : T100;
  assign T100 = T264 ? 8'h85 : T101;
  assign T101 = T263 ? 8'h86 : T102;
  assign T102 = T262 ? 8'h87 : T103;
  assign T103 = T261 ? 8'h88 : T104;
  assign T104 = T260 ? 8'h89 : T105;
  assign T105 = T259 ? 8'h8a : T106;
  assign T106 = T258 ? 8'h8b : T107;
  assign T107 = T257 ? 8'h8c : T108;
  assign T108 = T256 ? 8'h8d : T109;
  assign T109 = T255 ? 8'h8e : T110;
  assign T110 = T254 ? 8'h8f : T111;
  assign T111 = T253 ? 8'h90 : T112;
  assign T112 = T252 ? 8'h91 : T113;
  assign T113 = T251 ? 8'h92 : T114;
  assign T114 = T250 ? 8'h93 : T115;
  assign T115 = T249 ? 8'h94 : T116;
  assign T116 = T248 ? 8'h95 : T117;
  assign T117 = T247 ? 8'h96 : T118;
  assign T118 = T246 ? 8'h97 : T119;
  assign T119 = T245 ? 8'h98 : T120;
  assign T120 = T244 ? 8'h99 : T121;
  assign T121 = T243 ? 8'h9a : T122;
  assign T122 = T242 ? 8'h9b : T123;
  assign T123 = T241 ? 8'h9c : T124;
  assign T124 = T240 ? 8'h9d : T125;
  assign T125 = T239 ? 8'h9e : T126;
  assign T126 = T127 ? 8'h9f : 8'ha0;
  assign T127 = T128[1'h1:1'h1];
  assign T128 = T761 ^ T129;
  assign T129 = T130 << 1'h1;
  assign T130 = 108'h0 | T131;
  assign T131 = sigSum[7'h6c:1'h1];
  assign sigSum = T760 + alignedNegSigC;
  assign alignedNegSigC = T132[8'ha1:1'h0];
  assign T132 = {T228, T133};
  assign T133 = T138 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T135 ^ T134;
  assign T134 = io_op[1'h0:1'h0];
  assign T135 = io_c[7'h40:7'h40];
  assign signProd = T137 ^ T136;
  assign T136 = io_op[1'h1:1'h1];
  assign T137 = signA ^ signB;
  assign signB = io_b[7'h40:7'h40];
  assign signA = io_a[7'h40:7'h40];
  assign T138 = T139 != 53'h0;
  assign T139 = sigC & CExtraMask;
  assign CExtraMask = {T195, T140};
  assign T140 = {T170, T141};
  assign T141 = {T160, T142};
  assign T142 = T143[3'h4:3'h4];
  assign T143 = T144[5'h14:5'h10];
  assign T144 = T145[6'h34:6'h20];
  assign T145 = T146[8'h93:7'h5f];
  assign T146 = $signed(257'h10000000000000000000000000000000000000000000000000000000000000000) >>> CAlignDist;
  assign CAlignDist = T147[3'h7:1'h0];
  assign T147 = CAlignDist_floor ? 14'h0 : T148;
  assign T148 = T155 ? sNatCAlignDist : 14'ha1;
  assign sNatCAlignDist = sExpAlignedProd - T747;
  assign T747 = {2'h0, expC};
  assign expC = io_c[6'h3f:6'h34];
  assign sExpAlignedProd = T149 + 14'h38;
  assign T149 = T150 + T748;
  assign T748 = {2'h0, expA};
  assign expA = io_a[6'h3f:6'h34];
  assign T150 = {T152, T151};
  assign T151 = expB[4'ha:1'h0];
  assign expB = io_b[6'h3f:6'h34];
  assign T152 = 3'h0 - T749;
  assign T749 = {2'h0, T153};
  assign T153 = T154 ^ 1'h1;
  assign T154 = expB[4'hb:4'hb];
  assign T155 = T156 < 13'ha1;
  assign T156 = sNatCAlignDist[4'hc:1'h0];
  assign CAlignDist_floor = isZeroProd | T157;
  assign T157 = sNatCAlignDist[4'hd:4'hd];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T158 == 3'h0;
  assign T158 = expB[4'hb:4'h9];
  assign isZeroA = T159 == 3'h0;
  assign T159 = expA[4'hb:4'h9];
  assign T160 = {T166, T161};
  assign T161 = {T165, T162};
  assign T162 = T163[1'h1:1'h1];
  assign T163 = T164[2'h3:2'h2];
  assign T164 = T143[2'h3:1'h0];
  assign T165 = T163[1'h0:1'h0];
  assign T166 = {T169, T167};
  assign T167 = T168[1'h1:1'h1];
  assign T168 = T164[1'h1:1'h0];
  assign T169 = T168[1'h0:1'h0];
  assign T170 = T193 | T171;
  assign T171 = T172 & 16'haaaa;
  assign T172 = T173 << 1'h1;
  assign T173 = T174[4'he:1'h0];
  assign T174 = T191 | T175;
  assign T175 = T176 & 16'hcccc;
  assign T176 = T177 << 2'h2;
  assign T177 = T178[4'hd:1'h0];
  assign T178 = T189 | T179;
  assign T179 = T180 & 16'hf0f0;
  assign T180 = T181 << 3'h4;
  assign T181 = T182[4'hb:1'h0];
  assign T182 = T187 | T183;
  assign T183 = T184 & 16'hff00;
  assign T184 = T185 << 4'h8;
  assign T185 = T186[3'h7:1'h0];
  assign T186 = T144[4'hf:1'h0];
  assign T187 = T750 & 16'hff;
  assign T750 = {8'h0, T188};
  assign T188 = T186 >> 4'h8;
  assign T189 = T751 & 16'hf0f;
  assign T751 = {4'h0, T190};
  assign T190 = T182 >> 3'h4;
  assign T191 = T752 & 16'h3333;
  assign T752 = {2'h0, T192};
  assign T192 = T178 >> 2'h2;
  assign T193 = T753 & 16'h5555;
  assign T753 = {1'h0, T194};
  assign T194 = T174 >> 1'h1;
  assign T195 = T224 | T196;
  assign T196 = T197 & 32'haaaaaaaa;
  assign T197 = T198 << 1'h1;
  assign T198 = T199[5'h1e:1'h0];
  assign T199 = T222 | T200;
  assign T200 = T201 & 32'hcccccccc;
  assign T201 = T202 << 2'h2;
  assign T202 = T203[5'h1d:1'h0];
  assign T203 = T220 | T204;
  assign T204 = T205 & 32'hf0f0f0f0;
  assign T205 = T206 << 3'h4;
  assign T206 = T207[5'h1b:1'h0];
  assign T207 = T218 | T208;
  assign T208 = T209 & 32'hff00ff00;
  assign T209 = T210 << 4'h8;
  assign T210 = T211[5'h17:1'h0];
  assign T211 = T216 | T212;
  assign T212 = T213 & 32'hffff0000;
  assign T213 = T214 << 5'h10;
  assign T214 = T215[4'hf:1'h0];
  assign T215 = T145[5'h1f:1'h0];
  assign T216 = T754 & 32'hffff;
  assign T754 = {16'h0, T217};
  assign T217 = T215 >> 5'h10;
  assign T218 = T755 & 32'hff00ff;
  assign T755 = {8'h0, T219};
  assign T219 = T211 >> 4'h8;
  assign T220 = T756 & 32'hf0f0f0f;
  assign T756 = {4'h0, T221};
  assign T221 = T207 >> 3'h4;
  assign T222 = T757 & 32'h33333333;
  assign T757 = {2'h0, T223};
  assign T223 = T203 >> 2'h2;
  assign T224 = T758 & 32'h55555555;
  assign T758 = {1'h0, T225};
  assign T225 = T199 >> 1'h1;
  assign sigC = {T226, fractC};
  assign fractC = io_c[6'h33:1'h0];
  assign T226 = isZeroC ^ 1'h1;
  assign isZeroC = T227 == 3'h0;
  assign T227 = expC[4'hb:4'h9];
  assign T228 = $signed(T229) >>> CAlignDist;
  assign T229 = T230;
  assign T230 = {doSubMags, T231};
  assign T231 = {negSigC, T232};
  assign T232 = 108'h0 - T759;
  assign T759 = {107'h0, doSubMags};
  assign negSigC = doSubMags ? T233 : sigC;
  assign T233 = ~ sigC;
  assign T760 = {55'h0, T234};
  assign T234 = T235 << 1'h1;
  assign T235 = sigA * sigB;
  assign sigB = {T236, fractB};
  assign fractB = io_b[6'h33:1'h0];
  assign T236 = isZeroB ^ 1'h1;
  assign sigA = {T237, fractA};
  assign fractA = io_a[6'h33:1'h0];
  assign T237 = isZeroA ^ 1'h1;
  assign T761 = {1'h0, T238};
  assign T238 = 108'h0 ^ T131;
  assign T239 = T128[2'h2:2'h2];
  assign T240 = T128[2'h3:2'h3];
  assign T241 = T128[3'h4:3'h4];
  assign T242 = T128[3'h5:3'h5];
  assign T243 = T128[3'h6:3'h6];
  assign T244 = T128[3'h7:3'h7];
  assign T245 = T128[4'h8:4'h8];
  assign T246 = T128[4'h9:4'h9];
  assign T247 = T128[4'ha:4'ha];
  assign T248 = T128[4'hb:4'hb];
  assign T249 = T128[4'hc:4'hc];
  assign T250 = T128[4'hd:4'hd];
  assign T251 = T128[4'he:4'he];
  assign T252 = T128[4'hf:4'hf];
  assign T253 = T128[5'h10:5'h10];
  assign T254 = T128[5'h11:5'h11];
  assign T255 = T128[5'h12:5'h12];
  assign T256 = T128[5'h13:5'h13];
  assign T257 = T128[5'h14:5'h14];
  assign T258 = T128[5'h15:5'h15];
  assign T259 = T128[5'h16:5'h16];
  assign T260 = T128[5'h17:5'h17];
  assign T261 = T128[5'h18:5'h18];
  assign T262 = T128[5'h19:5'h19];
  assign T263 = T128[5'h1a:5'h1a];
  assign T264 = T128[5'h1b:5'h1b];
  assign T265 = T128[5'h1c:5'h1c];
  assign T266 = T128[5'h1d:5'h1d];
  assign T267 = T128[5'h1e:5'h1e];
  assign T268 = T128[5'h1f:5'h1f];
  assign T269 = T128[6'h20:6'h20];
  assign T270 = T128[6'h21:6'h21];
  assign T271 = T128[6'h22:6'h22];
  assign T272 = T128[6'h23:6'h23];
  assign T273 = T128[6'h24:6'h24];
  assign T274 = T128[6'h25:6'h25];
  assign T275 = T128[6'h26:6'h26];
  assign T276 = T128[6'h27:6'h27];
  assign T277 = T128[6'h28:6'h28];
  assign T278 = T128[6'h29:6'h29];
  assign T279 = T128[6'h2a:6'h2a];
  assign T280 = T128[6'h2b:6'h2b];
  assign T281 = T128[6'h2c:6'h2c];
  assign T282 = T128[6'h2d:6'h2d];
  assign T283 = T128[6'h2e:6'h2e];
  assign T284 = T128[6'h2f:6'h2f];
  assign T285 = T128[6'h30:6'h30];
  assign T286 = T128[6'h31:6'h31];
  assign T287 = T128[6'h32:6'h32];
  assign T288 = T128[6'h33:6'h33];
  assign T289 = T128[6'h34:6'h34];
  assign T290 = T128[6'h35:6'h35];
  assign T291 = T128[6'h36:6'h36];
  assign T292 = T128[6'h37:6'h37];
  assign T293 = T128[6'h38:6'h38];
  assign T294 = T128[6'h39:6'h39];
  assign T295 = T128[6'h3a:6'h3a];
  assign T296 = T128[6'h3b:6'h3b];
  assign T297 = T128[6'h3c:6'h3c];
  assign T298 = T128[6'h3d:6'h3d];
  assign T299 = T128[6'h3e:6'h3e];
  assign T300 = T128[6'h3f:6'h3f];
  assign T301 = T128[7'h40:7'h40];
  assign T302 = T128[7'h41:7'h41];
  assign T303 = T128[7'h42:7'h42];
  assign T304 = T128[7'h43:7'h43];
  assign T305 = T128[7'h44:7'h44];
  assign T306 = T128[7'h45:7'h45];
  assign T307 = T128[7'h46:7'h46];
  assign T308 = T128[7'h47:7'h47];
  assign T309 = T128[7'h48:7'h48];
  assign T310 = T128[7'h49:7'h49];
  assign T311 = T128[7'h4a:7'h4a];
  assign T312 = T128[7'h4b:7'h4b];
  assign T313 = T128[7'h4c:7'h4c];
  assign T314 = T128[7'h4d:7'h4d];
  assign T315 = T128[7'h4e:7'h4e];
  assign T316 = T128[7'h4f:7'h4f];
  assign T317 = T128[7'h50:7'h50];
  assign T318 = T128[7'h51:7'h51];
  assign T319 = T128[7'h52:7'h52];
  assign T320 = T128[7'h53:7'h53];
  assign T321 = T128[7'h54:7'h54];
  assign T322 = T128[7'h55:7'h55];
  assign T323 = T128[7'h56:7'h56];
  assign T324 = T128[7'h57:7'h57];
  assign T325 = T128[7'h58:7'h58];
  assign T326 = T128[7'h59:7'h59];
  assign T327 = T128[7'h5a:7'h5a];
  assign T328 = T128[7'h5b:7'h5b];
  assign T329 = T128[7'h5c:7'h5c];
  assign T330 = T128[7'h5d:7'h5d];
  assign T331 = T128[7'h5e:7'h5e];
  assign T332 = T128[7'h5f:7'h5f];
  assign T333 = T128[7'h60:7'h60];
  assign T334 = T128[7'h61:7'h61];
  assign T335 = T128[7'h62:7'h62];
  assign T336 = T128[7'h63:7'h63];
  assign T337 = T128[7'h64:7'h64];
  assign T338 = T128[7'h65:7'h65];
  assign T339 = T128[7'h66:7'h66];
  assign T340 = T128[7'h67:7'h67];
  assign T341 = T128[7'h68:7'h68];
  assign T342 = T128[7'h69:7'h69];
  assign T343 = T128[7'h6a:7'h6a];
  assign T344 = T128[7'h6b:7'h6b];
  assign notCDom_signSigSum = sigSum[7'h6d:7'h6d];
  assign CDom_estNormDist = T347 ? CAlignDist : T762;
  assign T762 = {2'h0, T345};
  assign T345 = T346[3'h5:1'h0];
  assign T346 = CAlignDist - 8'h1;
  assign T347 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T348;
  assign T348 = T349 == 13'h0;
  assign T349 = sNatCAlignDist[4'hc:1'h0];
  assign isCDominant = T353 & T350;
  assign T350 = CAlignDist_floor | T351;
  assign T351 = T352 < 13'h36;
  assign T352 = sNatCAlignDist[4'hc:1'h0];
  assign T353 = isZeroC ^ 1'h1;
  assign sExpSum = CAlignDist_floor ? T763 : sExpAlignedProd;
  assign T763 = {2'h0, expC};
  assign T354 = T14[1'h0:1'h0];
  assign T355 = {T361, T356};
  assign T356 = {T360, T357};
  assign T357 = T358[1'h1:1'h1];
  assign T358 = T359[2'h3:2'h2];
  assign T359 = T15[2'h3:1'h0];
  assign T360 = T358[1'h0:1'h0];
  assign T361 = {T364, T362};
  assign T362 = T363[1'h1:1'h1];
  assign T363 = T359[1'h1:1'h0];
  assign T364 = T363[1'h0:1'h0];
  assign T365 = T388 | T366;
  assign T366 = T367 & 16'haaaa;
  assign T367 = T368 << 1'h1;
  assign T368 = T369[4'he:1'h0];
  assign T369 = T386 | T370;
  assign T370 = T371 & 16'hcccc;
  assign T371 = T372 << 2'h2;
  assign T372 = T373[4'hd:1'h0];
  assign T373 = T384 | T374;
  assign T374 = T375 & 16'hf0f0;
  assign T375 = T376 << 3'h4;
  assign T376 = T377[4'hb:1'h0];
  assign T377 = T382 | T378;
  assign T378 = T379 & 16'hff00;
  assign T379 = T380 << 4'h8;
  assign T380 = T381[3'h7:1'h0];
  assign T381 = T16[4'hf:1'h0];
  assign T382 = T764 & 16'hff;
  assign T764 = {8'h0, T383};
  assign T383 = T381 >> 4'h8;
  assign T384 = T765 & 16'hf0f;
  assign T765 = {4'h0, T385};
  assign T385 = T377 >> 3'h4;
  assign T386 = T766 & 16'h3333;
  assign T766 = {2'h0, T387};
  assign T387 = T373 >> 2'h2;
  assign T388 = T767 & 16'h5555;
  assign T767 = {1'h0, T389};
  assign T389 = T369 >> 1'h1;
  assign T390 = T419 | T391;
  assign T391 = T392 & 32'haaaaaaaa;
  assign T392 = T393 << 1'h1;
  assign T393 = T394[5'h1e:1'h0];
  assign T394 = T417 | T395;
  assign T395 = T396 & 32'hcccccccc;
  assign T396 = T397 << 2'h2;
  assign T397 = T398[5'h1d:1'h0];
  assign T398 = T415 | T399;
  assign T399 = T400 & 32'hf0f0f0f0;
  assign T400 = T401 << 3'h4;
  assign T401 = T402[5'h1b:1'h0];
  assign T402 = T413 | T403;
  assign T403 = T404 & 32'hff00ff00;
  assign T404 = T405 << 4'h8;
  assign T405 = T406[5'h17:1'h0];
  assign T406 = T411 | T407;
  assign T407 = T408 & 32'hffff0000;
  assign T408 = T409 << 5'h10;
  assign T409 = T410[4'hf:1'h0];
  assign T410 = T17[5'h1f:1'h0];
  assign T411 = T768 & 32'hffff;
  assign T768 = {16'h0, T412};
  assign T412 = T410 >> 5'h10;
  assign T413 = T769 & 32'hff00ff;
  assign T769 = {8'h0, T414};
  assign T414 = T406 >> 4'h8;
  assign T415 = T770 & 32'hf0f0f0f;
  assign T770 = {4'h0, T416};
  assign T416 = T402 >> 3'h4;
  assign T417 = T771 & 32'h33333333;
  assign T771 = {2'h0, T418};
  assign T418 = T398 >> 2'h2;
  assign T419 = T772 & 32'h55555555;
  assign T772 = {1'h0, T420};
  assign T420 = T394 >> 1'h1;
  assign T421 = 56'h0 - T773;
  assign T773 = {55'h0, T422};
  assign T422 = sExpX3[4'hd:4'hd];
  assign sigX3 = T423[6'h38:1'h0];
  assign T423 = {T595, T424};
  assign T424 = doIncrSig ? T591 : T425;
  assign T425 = T426 != 32'h0;
  assign T426 = T496 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T427, 1'h1};
  assign T427 = {T471, T428};
  assign T428 = {T452, T429};
  assign T429 = {T442, T430};
  assign T430 = {T438, T431};
  assign T431 = T432[2'h2:2'h2];
  assign T432 = T433[3'h6:3'h4];
  assign T433 = T434[4'he:4'h8];
  assign T434 = T435[5'h1e:5'h10];
  assign T435 = T436[5'h1f:1'h1];
  assign T436 = $signed(33'h100000000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T437;
  assign T437 = estNormDist[3'h4:1'h0];
  assign T438 = {T441, T439};
  assign T439 = T440[1'h1:1'h1];
  assign T440 = T432[1'h1:1'h0];
  assign T441 = T440[1'h0:1'h0];
  assign T442 = {T448, T443};
  assign T443 = {T447, T444};
  assign T444 = T445[1'h1:1'h1];
  assign T445 = T446[2'h3:2'h2];
  assign T446 = T433[2'h3:1'h0];
  assign T447 = T445[1'h0:1'h0];
  assign T448 = {T451, T449};
  assign T449 = T450[1'h1:1'h1];
  assign T450 = T446[1'h1:1'h0];
  assign T451 = T450[1'h0:1'h0];
  assign T452 = T469 | T453;
  assign T453 = T454 & 8'haa;
  assign T454 = T455 << 1'h1;
  assign T455 = T456[3'h6:1'h0];
  assign T456 = T467 | T457;
  assign T457 = T458 & 8'hcc;
  assign T458 = T459 << 2'h2;
  assign T459 = T460[3'h5:1'h0];
  assign T460 = T465 | T461;
  assign T461 = T462 & 8'hf0;
  assign T462 = T463 << 3'h4;
  assign T463 = T464[2'h3:1'h0];
  assign T464 = T434[3'h7:1'h0];
  assign T465 = T774 & 8'hf;
  assign T774 = {4'h0, T466};
  assign T466 = T464 >> 3'h4;
  assign T467 = T775 & 8'h33;
  assign T775 = {2'h0, T468};
  assign T468 = T460 >> 2'h2;
  assign T469 = T776 & 8'h55;
  assign T776 = {1'h0, T470};
  assign T470 = T456 >> 1'h1;
  assign T471 = T494 | T472;
  assign T472 = T473 & 16'haaaa;
  assign T473 = T474 << 1'h1;
  assign T474 = T475[4'he:1'h0];
  assign T475 = T492 | T476;
  assign T476 = T477 & 16'hcccc;
  assign T477 = T478 << 2'h2;
  assign T478 = T479[4'hd:1'h0];
  assign T479 = T490 | T480;
  assign T480 = T481 & 16'hf0f0;
  assign T481 = T482 << 3'h4;
  assign T482 = T483[4'hb:1'h0];
  assign T483 = T488 | T484;
  assign T484 = T485 & 16'hff00;
  assign T485 = T486 << 4'h8;
  assign T486 = T487[3'h7:1'h0];
  assign T487 = T435[4'hf:1'h0];
  assign T488 = T777 & 16'hff;
  assign T777 = {8'h0, T489};
  assign T489 = T487 >> 4'h8;
  assign T490 = T778 & 16'hf0f;
  assign T778 = {4'h0, T491};
  assign T491 = T483 >> 3'h4;
  assign T492 = T779 & 16'h3333;
  assign T779 = {2'h0, T493};
  assign T493 = T479 >> 2'h2;
  assign T494 = T780 & 16'h5555;
  assign T780 = {1'h0, T495};
  assign T495 = T475 >> 1'h1;
  assign T496 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T570 : T781;
  assign T781 = {1'h0, T497};
  assign T497 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T534 ? T522 : T498;
  assign T498 = T521 ? T502 : T499;
  assign T499 = {T501, T500};
  assign T500 = 54'h0 - T782;
  assign T782 = {53'h0, doSubMags};
  assign T501 = sigSum[6'h21:1'h1];
  assign T502 = T520 ? T784 : T503;
  assign T503 = {T505, T504};
  assign T504 = 86'h0 - T783;
  assign T783 = {85'h0, doSubMags};
  assign T505 = sigSum[1'h1:1'h1];
  assign T784 = {21'h0, T506};
  assign T506 = {T519, T507};
  assign T507 = doSubMags ? T513 : T508;
  assign T508 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T511, T509};
  assign T509 = T510 != 44'h0;
  assign T510 = sigSum[6'h2b:1'h0];
  assign T511 = T512 != 32'h0;
  assign T512 = sigSum[7'h4b:6'h2c];
  assign T513 = ~ T514;
  assign T514 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T517, T515};
  assign T515 = T516 != 44'h0;
  assign T516 = notSigSum[6'h2b:1'h0];
  assign notSigSum = ~ sigSum;
  assign T517 = T518 != 32'h0;
  assign T518 = notSigSum[7'h4b:6'h2c];
  assign T519 = sigSum[7'h6c:6'h2c];
  assign T520 = estNormNeg_dist[3'h4:3'h4];
  assign T521 = estNormNeg_dist[3'h5:3'h5];
  assign T522 = T533 ? T530 : T523;
  assign T523 = {T529, T524};
  assign T524 = doSubMags ? T527 : T525;
  assign T525 = T526 != 11'h0;
  assign T526 = sigSum[4'hb:1'h1];
  assign T527 = T528 == 11'h0;
  assign T528 = notSigSum[4'hb:1'h1];
  assign T529 = sigSum[7'h61:4'hc];
  assign T530 = {T532, T531};
  assign T531 = 22'h0 - T785;
  assign T785 = {21'h0, doSubMags};
  assign T532 = sigSum[7'h41:1'h1];
  assign T533 = estNormNeg_dist[3'h5:3'h5];
  assign T534 = estNormNeg_dist[3'h6:3'h6];
  assign CDom_firstNormAbsSigSum = T535;
  assign T535 = T543 | T536;
  assign T536 = T786 & T537;
  assign T537 = {T539, T538};
  assign T538 = firstReduceNotSigSum[1'h0:1'h0];
  assign T539 = notSigSum[8'h81:6'h2c];
  assign T786 = T540 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T540 = T541;
  assign T541 = doSubMags & T542;
  assign T542 = CDom_estNormDist[3'h5:3'h5];
  assign T543 = T552 | T544;
  assign T544 = T787 & T545;
  assign T545 = {T547, T546};
  assign T546 = firstReduceNotSigSum != 2'h0;
  assign T547 = notSigSum[8'ha1:7'h4c];
  assign T787 = T548 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T548 = T549;
  assign T549 = doSubMags & T550;
  assign T550 = ~ T551;
  assign T551 = CDom_estNormDist[3'h5:3'h5];
  assign T552 = T561 | T553;
  assign T553 = T788 & T554;
  assign T554 = {T556, T555};
  assign T555 = firstReduceSigSum[1'h0:1'h0];
  assign T556 = sigSum[8'h81:6'h2c];
  assign T788 = T557 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T557 = T558;
  assign T558 = T560 & T559;
  assign T559 = CDom_estNormDist[3'h5:3'h5];
  assign T560 = ~ doSubMags;
  assign T561 = T789 & T562;
  assign T562 = {T564, T563};
  assign T563 = firstReduceSigSum != 2'h0;
  assign T564 = sigSum[8'ha1:7'h4c];
  assign T789 = T565 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T565 = T566;
  assign T566 = T569 & T567;
  assign T567 = ~ T568;
  assign T568 = CDom_estNormDist[3'h5:3'h5];
  assign T569 = ~ doSubMags;
  assign T570 = isCDominant ? T791 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T590 ? T582 : T571;
  assign T571 = T581 ? T574 : T572;
  assign T572 = T573 << 6'h36;
  assign T573 = notSigSum[6'h22:1'h1];
  assign T574 = T580 ? T790 : T575;
  assign T575 = T576 << 7'h56;
  assign T576 = notSigSum[2'h2:1'h1];
  assign T790 = {23'h0, T577};
  assign T577 = {T579, T578};
  assign T578 = firstReduceNotSigSum[1'h0:1'h0];
  assign T579 = notSigSum[7'h6b:6'h2c];
  assign T580 = estNormNeg_dist[3'h4:3'h4];
  assign T581 = estNormNeg_dist[3'h5:3'h5];
  assign T582 = T589 ? T587 : T583;
  assign T583 = {T586, T584};
  assign T584 = T585 != 11'h0;
  assign T585 = notSigSum[4'hb:1'h1];
  assign T586 = notSigSum[7'h62:4'hc];
  assign T587 = T588 << 5'h16;
  assign T588 = notSigSum[7'h42:1'h1];
  assign T589 = estNormNeg_dist[3'h5:3'h5];
  assign T590 = estNormNeg_dist[3'h6:3'h6];
  assign T791 = {1'h0, CDom_firstNormAbsSigSum};
  assign T591 = T592 == 32'h0;
  assign T592 = T593 & absSigSumExtraMask;
  assign T593 = ~ T594;
  assign T594 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign T595 = T596 >> normTo2ShiftDist;
  assign T596 = cFirstNormAbsSigSum[7'h57:1'h1];
  assign roundPosBit = T597 != 57'h0;
  assign T597 = sigX3 & T792;
  assign T792 = {1'h0, roundPosMask};
  assign roundPosMask = T793 & roundMask;
  assign T793 = {1'h0, T598};
  assign T598 = ~ T599;
  assign T599 = roundMask >> 1'h1;
  assign T600 = ~ allRound;
  assign allRound = roundPosBit & allRoundExtra;
  assign allRoundExtra = T601 == 57'h0;
  assign T601 = T603 & T794;
  assign T794 = {2'h0, T602};
  assign T602 = roundMask >> 1'h1;
  assign T603 = ~ sigX3;
  assign doIncrSig = T604 & doSubMags;
  assign T604 = T606 & T605;
  assign T605 = ~ notCDom_signSigSum;
  assign T606 = ~ isCDominant;
  assign commonCase = T608 & T607;
  assign T607 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T608 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T609 == 2'h3;
  assign T609 = expC[4'hb:4'ha];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T610 == 2'h3;
  assign T610 = expB[4'hb:4'ha];
  assign isSpecialA = T611 == 2'h3;
  assign T611 = expA[4'hb:4'ha];
  assign underflow = commonCase & underflowY;
  assign underflowY = inexactY & T612;
  assign T612 = T616 | T613;
  assign T613 = sExpX3_13 <= T795;
  assign T795 = {2'h0, T614};
  assign T614 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign sigX3Shift1 = T615 == 2'h0;
  assign T615 = sigX3[6'h38:6'h37];
  assign T616 = sExpX3[4'hd:4'hd];
  assign overflow = commonCase & overflowY;
  assign overflowY = T617 == 3'h3;
  assign T617 = sExpY[4'hc:4'ha];
  assign sExpY = T664 | T618;
  assign T618 = T620 ? T619 : 14'h0;
  assign T619 = sExpX3 - 14'h1;
  assign T620 = T621 == 2'h0;
  assign T621 = sigY3[6'h36:6'h35];
  assign sigY3 = T635 | T622;
  assign T622 = roundEven ? T623 : 55'h0;
  assign T623 = roundUp_sigY3 & T624;
  assign T624 = ~ T625;
  assign T625 = roundMask >> 1'h1;
  assign roundUp_sigY3 = T626[6'h36:1'h0];
  assign T626 = T627 + 55'h1;
  assign T627 = T628 >> 2'h2;
  assign T628 = sigX3 | T796;
  assign T796 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T632 : T629;
  assign T629 = T631 & T630;
  assign T630 = ~ anyRoundExtra;
  assign T631 = roundingMode_nearest_even & roundPosBit;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T632 = T633 & allRoundExtra;
  assign T633 = roundingMode_nearest_even & T634;
  assign T634 = ~ roundPosBit;
  assign T635 = T657 | T636;
  assign T636 = roundUp ? roundUp_sigY3 : 55'h0;
  assign roundUp = T644 | T637;
  assign T637 = T638 & 1'h1;
  assign T638 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T642 & T639;
  assign T639 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T640 : notCDom_signSigSum;
  assign T640 = doSubMags & T641;
  assign T641 = ~ isZeroC;
  assign T642 = ~ isZeroY;
  assign isZeroY = T643 == 3'h0;
  assign T643 = sigX3[6'h38:6'h36];
  assign T644 = T647 | T645;
  assign T645 = T646 & roundPosBit;
  assign T646 = doIncrSig & roundingMode_nearest_even;
  assign T647 = T649 | T648;
  assign T648 = doIncrSig & allRound;
  assign T649 = T653 | T650;
  assign T650 = T651 & anyRound;
  assign T651 = T652 & roundDirectUp;
  assign T652 = ~ doIncrSig;
  assign T653 = T654 & anyRoundExtra;
  assign T654 = T655 & roundPosBit;
  assign T655 = T656 & roundingMode_nearest_even;
  assign T656 = ~ doIncrSig;
  assign T657 = T661 ? T658 : 55'h0;
  assign T658 = T659 >> 2'h2;
  assign T659 = sigX3 & T797;
  assign T797 = {1'h0, T660};
  assign T660 = ~ roundMask;
  assign T661 = T663 & T662;
  assign T662 = ~ roundEven;
  assign T663 = ~ roundUp;
  assign T664 = T667 | T665;
  assign T665 = T666 ? sExpX3 : 14'h0;
  assign T666 = sigY3[6'h35:6'h35];
  assign T667 = T669 ? T668 : 14'h0;
  assign T668 = sExpX3 + 14'h1;
  assign T669 = sigY3[6'h36:6'h36];
  assign T670 = {invalid, 1'h0};
  assign invalid = T689 | notSigNaN_invalid;
  assign notSigNaN_invalid = T686 | T671;
  assign T671 = T672 & doSubMags;
  assign T672 = T675 & isInfC;
  assign isInfC = isSpecialC & T673;
  assign T673 = T674 ^ 1'h1;
  assign T674 = expC[4'h9:4'h9];
  assign T675 = T681 & T676;
  assign T676 = isInfA | isInfB;
  assign isInfB = isSpecialB & T677;
  assign T677 = T678 ^ 1'h1;
  assign T678 = expB[4'h9:4'h9];
  assign isInfA = isSpecialA & T679;
  assign T679 = T680 ^ 1'h1;
  assign T680 = expA[4'h9:4'h9];
  assign T681 = T684 & T682;
  assign T682 = ~ isNaNB;
  assign isNaNB = isSpecialB & T683;
  assign T683 = expB[4'h9:4'h9];
  assign T684 = ~ isNaNA;
  assign isNaNA = isSpecialA & T685;
  assign T685 = expA[4'h9:4'h9];
  assign T686 = T688 | T687;
  assign T687 = isZeroA & isInfB;
  assign T688 = isInfA & isZeroB;
  assign T689 = T693 | isSigNaNC;
  assign isSigNaNC = isNaNC & T690;
  assign T690 = T691 ^ 1'h1;
  assign T691 = fractC[6'h33:6'h33];
  assign isNaNC = isSpecialC & T692;
  assign T692 = expC[4'h9:4'h9];
  assign T693 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T694;
  assign T694 = T695 ^ 1'h1;
  assign T695 = fractB[6'h33:6'h33];
  assign isSigNaNA = isNaNA & T696;
  assign T696 = T697 ^ 1'h1;
  assign T697 = fractA[6'h33:6'h33];
  assign io_out = T698;
  assign T698 = {signOut, T699};
  assign T699 = {expOut, fractOut};
  assign fractOut = fractY | T700;
  assign T700 = 52'h0 - T798;
  assign T798 = {51'h0, T701};
  assign T701 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T702;
  assign T702 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T705 | T703;
  assign T703 = roundingMode_max & T704;
  assign T704 = ~ signY;
  assign T705 = roundingMode_nearest_even | T706;
  assign T706 = roundingMode_min & signY;
  assign isNaNOut = T707 | notSigNaN_invalid;
  assign T707 = T708 | isNaNC;
  assign T708 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T710 : T709;
  assign T709 = sigY3[6'h34:1'h1];
  assign T710 = sigY3[6'h33:1'h0];
  assign expOut = T712 | T711;
  assign T711 = isNaNOut ? 12'he00 : 12'h0;
  assign T712 = T717 | T713;
  assign T713 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = T715 | T714;
  assign T714 = overflow & overflowY_roundMagUp;
  assign T715 = T716 | isInfC;
  assign T716 = isInfA | isInfB;
  assign T717 = T719 | T718;
  assign T718 = isSatOut ? 12'hbff : 12'h0;
  assign T719 = T722 & T720;
  assign T720 = ~ T721;
  assign T721 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T722 = T725 & T723;
  assign T723 = ~ T724;
  assign T724 = isSatOut ? 12'h400 : 12'h0;
  assign T725 = expY & T726;
  assign T726 = ~ T727;
  assign T727 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign notSpecial_isZeroOut = T731 | totalUnderflowY;
  assign totalUnderflowY = T730 | T728;
  assign T728 = T729 < 12'h3ce;
  assign T729 = sExpY[4'hb:1'h0];
  assign T730 = sExpY[4'hc:4'hc];
  assign T731 = notSpecial_addZeros | isZeroY;
  assign expY = sExpY[4'hb:1'h0];
  assign signOut = T733 | T732;
  assign T732 = commonCase & signY;
  assign T733 = T737 | T734;
  assign T734 = T735 & opSignC;
  assign T735 = T736 & isSpecialC;
  assign T736 = mulSpecial ^ 1'h1;
  assign T737 = T741 | T738;
  assign T738 = T739 & signProd;
  assign T739 = mulSpecial & T740;
  assign T740 = isSpecialC ^ 1'h1;
  assign T741 = T742 | isNaNOut;
  assign T742 = T743 & opSignC;
  assign T743 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_1(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T30;
  reg [2:0] in_rm;
  wire[2:0] T0;
  reg [64:0] in_in3;
  wire[64:0] T1;
  wire[64:0] T2;
  wire[64:0] zero;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg [64:0] in_in2;
  wire[64:0] T9;
  wire[64:0] T10;
  wire T11;
  reg [64:0] in_in1;
  wire[64:0] T12;
  wire[1:0] T31;
  reg [4:0] in_cmd;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[4:0] T32;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [4:0] R20;
  wire[4:0] T21;
  reg [4:0] R22;
  wire[4:0] T23;
  wire[4:0] res_exc;
  reg  valid;
  reg  R24;
  wire T33;
  reg [64:0] R25;
  wire[64:0] T26;
  reg [64:0] R27;
  wire[64:0] T28;
  wire[64:0] res_data;
  reg  R29;
  wire T34;
  wire[64:0] fma_io_out;
  wire[4:0] fma_io_exceptionFlags;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R20 = {1{$random}};
    R22 = {1{$random}};
    valid = {1{$random}};
    R24 = {1{$random}};
    R25 = {3{$random}};
    R27 = {3{$random}};
    R29 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T30 = in_rm[1'h1:1'h0];
  assign T0 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T1 = T6 ? zero : T2;
  assign T2 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign zero = T3 << 7'h40;
  assign T3 = T5 ^ T4;
  assign T4 = io_in_bits_in2[7'h40:7'h40];
  assign T5 = io_in_bits_in1[7'h40:7'h40];
  assign T6 = io_in_valid & T7;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T9 = T11 ? 65'h8000000000000000 : T10;
  assign T10 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T11 = io_in_valid & io_in_bits_swap23;
  assign T12 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T31 = in_cmd[1'h1:1'h0];
  assign T13 = io_in_valid ? T32 : T14;
  assign T14 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T32 = {3'h0, T15};
  assign T15 = {T17, T16};
  assign T16 = io_in_bits_cmd[1'h0:1'h0];
  assign T17 = T19 & T18;
  assign T18 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T19 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R20;
  assign T21 = R24 ? R22 : R20;
  assign T23 = valid ? res_exc : R22;
  assign res_exc = fma_io_exceptionFlags;
  assign T33 = reset ? 1'h0 : valid;
  assign io_out_bits_data = R25;
  assign T26 = R24 ? R27 : R25;
  assign T28 = valid ? res_data : R27;
  assign res_data = fma_io_out;
  assign io_out_valid = R29;
  assign T34 = reset ? 1'h0 : R24;
  mulAddSubRecodedFloatN_1 fma(
       .io_op( T31 ),
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_c( in_in3 ),
       .io_roundingMode( T30 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T6) begin
      in_in3 <= zero;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T11) begin
      in_in2 <= 65'h8000000000000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T32;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(R24) begin
      R20 <= R22;
    end
    if(valid) begin
      R22 <= res_exc;
    end
    valid <= io_in_valid;
    if(reset) begin
      R24 <= 1'h0;
    end else begin
      R24 <= valid;
    end
    if(R24) begin
      R25 <= R27;
    end
    if(valid) begin
      R27 <= res_data;
    end
    if(reset) begin
      R29 <= 1'h0;
    end else begin
      R29 <= R24;
    end
  end
endmodule

module recodedFloatNCompare(
    input [64:0] io_a,
    input [64:0] io_b,
    output io_a_eq_b,
    output io_a_lt_b,
    output io_a_eq_b_invalid,
    output io_a_lt_b_invalid
);

  wire T0;
  wire isNaNB;
  wire[2:0] codeB;
  wire[11:0] expB;
  wire isNaNA;
  wire[2:0] codeA;
  wire[11:0] expA;
  wire T1;
  wire isSignalingNaNB;
  wire T2;
  wire T3;
  wire[51:0] sigB;
  wire isSignalingNaNA;
  wire T4;
  wire T5;
  wire[51:0] sigA;
  wire T6;
  wire T7;
  wire T8;
  wire magLess;
  wire T9;
  wire T10;
  wire expEqual;
  wire T11;
  wire T12;
  wire T13;
  wire isZeroB;
  wire T14;
  wire isZeroA;
  wire T15;
  wire signA;
  wire T16;
  wire T17;
  wire magEqual;
  wire T18;
  wire T19;
  wire T20;
  wire signB;
  wire T21;
  wire T22;
  wire T23;
  wire signEqual;
  wire T24;
  wire T25;


  assign io_a_lt_b_invalid = T0;
  assign T0 = isNaNA | isNaNB;
  assign isNaNB = codeB == 3'h7;
  assign codeB = expB[4'hb:4'h9];
  assign expB = io_b[6'h3f:6'h34];
  assign isNaNA = codeA == 3'h7;
  assign codeA = expA[4'hb:4'h9];
  assign expA = io_a[6'h3f:6'h34];
  assign io_a_eq_b_invalid = T1;
  assign T1 = isSignalingNaNA | isSignalingNaNB;
  assign isSignalingNaNB = isNaNB & T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = sigB[6'h33:6'h33];
  assign sigB = io_b[6'h33:1'h0];
  assign isSignalingNaNA = isNaNA & T4;
  assign T4 = T5 ^ 1'h1;
  assign T5 = sigA[6'h33:6'h33];
  assign sigA = io_a[6'h33:1'h0];
  assign io_a_lt_b = T6;
  assign T6 = T21 & T7;
  assign T7 = signB ? T16 : T8;
  assign T8 = signA ? T12 : magLess;
  assign magLess = T11 | T9;
  assign T9 = expEqual & T10;
  assign T10 = sigA < sigB;
  assign expEqual = expA == expB;
  assign T11 = expA < expB;
  assign T12 = T13 ^ 1'h1;
  assign T13 = isZeroA & isZeroB;
  assign isZeroB = T14 ^ 1'h1;
  assign T14 = codeB != 3'h0;
  assign isZeroA = T15 ^ 1'h1;
  assign T15 = codeA != 3'h0;
  assign signA = io_a[7'h40:7'h40];
  assign T16 = T19 & T17;
  assign T17 = magEqual ^ 1'h1;
  assign magEqual = expEqual & T18;
  assign T18 = sigA == sigB;
  assign T19 = signA & T20;
  assign T20 = magLess ^ 1'h1;
  assign signB = io_b[7'h40:7'h40];
  assign T21 = io_a_lt_b_invalid ^ 1'h1;
  assign io_a_eq_b = T22;
  assign T22 = T24 & T23;
  assign T23 = isZeroA | signEqual;
  assign signEqual = signA == signB;
  assign T24 = T25 & magEqual;
  assign T25 = isNaNA ^ 1'h1;
endmodule

module FPToInt(input clk,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output io_out_bits_lt,
    output[63:0] io_out_bits_store,
    output[63:0] io_out_bits_toint,
    output[4:0] io_out_bits_exc
);

  reg [64:0] in_in2;
  wire[64:0] T0;
  wire[64:0] T1;
  wire[64:0] T2;
  wire[63:0] T3;
  wire[51:0] T4;
  wire[51:0] T5;
  wire[22:0] T6;
  wire[51:0] T7;
  wire[51:0] T352;
  wire T8;
  wire[2:0] T9;
  wire[11:0] T10;
  wire[11:0] T11;
  wire[11:0] T12;
  wire[11:0] T13;
  wire T14;
  wire[11:0] T15;
  wire[7:0] T19;
  wire T16;
  wire[11:0] T353;
  wire[10:0] T17;
  wire T18;
  wire[11:0] T354;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[4:0] T26;
  wire T27;
  wire T28;
  reg [64:0] in_in1;
  wire[64:0] T29;
  wire[64:0] T30;
  wire[64:0] T31;
  wire[63:0] T32;
  wire[51:0] T33;
  wire[51:0] T34;
  wire[22:0] T35;
  wire[51:0] T36;
  wire[51:0] T355;
  wire T37;
  wire[2:0] T38;
  wire[11:0] T39;
  wire[11:0] T40;
  wire[11:0] T41;
  wire[11:0] T42;
  wire T43;
  wire[11:0] T44;
  wire[7:0] T48;
  wire T45;
  wire[11:0] T356;
  wire[10:0] T46;
  wire T47;
  wire[11:0] T357;
  wire T49;
  wire T50;
  wire[4:0] T51;
  wire[4:0] T52;
  wire[4:0] dcmp_exc;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T358;
  wire[1:0] T55;
  wire[2:0] T56;
  reg [2:0] in_rm;
  wire[2:0] T57;
  wire T58;
  wire[4:0] T59;
  reg [4:0] in_cmd;
  wire[4:0] T60;
  wire[4:0] T61;
  wire[3:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire[1:0] T66;
  wire[2:0] T67;
  wire T68;
  wire[50:0] T69;
  wire[115:0] T70;
  wire[5:0] T71;
  wire[5:0] T72;
  wire[11:0] T73;
  wire T74;
  wire T75;
  wire[52:0] T76;
  wire[51:0] T77;
  wire T78;
  wire[1:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire[10:0] T88;
  wire T89;
  wire T90;
  wire[63:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[2:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[1:0] T109;
  wire T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[10:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  reg [1:0] in_typ;
  wire[1:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire[1:0] T149;
  wire T150;
  wire[4:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[63:0] T154;
  wire[63:0] unrec_out;
  wire[63:0] unrec_d;
  wire[62:0] T155;
  wire[51:0] T156;
  wire[51:0] T157;
  wire[51:0] T158;
  wire[52:0] T159;
  wire[5:0] T160;
  wire[5:0] T161;
  wire[11:0] T162;
  wire[52:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire[9:0] T167;
  wire T168;
  wire[1:0] T169;
  wire T170;
  wire[2:0] T171;
  wire[51:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire[1:0] T177;
  wire T178;
  wire T179;
  wire[1:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[10:0] T185;
  wire[10:0] T186;
  wire[10:0] T359;
  wire[10:0] T187;
  wire[10:0] T188;
  wire T189;
  wire[63:0] T190;
  wire[31:0] unrec_s;
  wire[30:0] T191;
  wire[22:0] T192;
  wire[22:0] T193;
  wire[22:0] T194;
  wire[23:0] T195;
  wire[4:0] T196;
  wire[4:0] T197;
  wire[8:0] T198;
  wire[23:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[6:0] T203;
  wire T204;
  wire[1:0] T205;
  wire T206;
  wire[2:0] T207;
  wire[22:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[1:0] T213;
  wire T214;
  wire T215;
  wire[1:0] T216;
  wire T217;
  wire T218;
  wire T219;
  wire[1:0] T220;
  wire[7:0] T221;
  wire[7:0] T222;
  wire[7:0] T360;
  wire[7:0] T223;
  wire[7:0] T224;
  wire T225;
  wire[31:0] T226;
  wire[31:0] T361;
  wire T227;
  reg  in_single;
  wire T228;
  wire[63:0] T362;
  wire[9:0] classify_out;
  wire[9:0] classify_d;
  wire[4:0] T229;
  wire[2:0] T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[11:0] T237;
  wire T238;
  wire[1:0] T239;
  wire[2:0] T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[9:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire[1:0] T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire[4:0] T259;
  wire[2:0] T260;
  wire[1:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[1:0] T268;
  wire T269;
  wire T270;
  wire T271;
  wire[51:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire[9:0] classify_s;
  wire[4:0] T276;
  wire[2:0] T277;
  wire[1:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[8:0] T284;
  wire T285;
  wire[1:0] T286;
  wire[2:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[6:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[1:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire[4:0] T306;
  wire[2:0] T307;
  wire[1:0] T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire[1:0] T315;
  wire T316;
  wire T317;
  wire T318;
  wire[22:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[63:0] T363;
  wire dcmp_out;
  wire[2:0] T324;
  wire[2:0] T364;
  wire[1:0] T325;
  wire[2:0] T326;
  wire[63:0] T327;
  wire[63:0] T365;
  wire[31:0] T328;
  wire[31:0] T329;
  wire[31:0] T366;
  wire T367;
  wire[63:0] T330;
  wire[63:0] T331;
  wire[63:0] T332;
  wire[63:0] T333;
  wire[63:0] T334;
  wire[63:0] T335;
  wire T336;
  wire[63:0] T337;
  wire[63:0] T338;
  wire[63:0] T339;
  wire[63:0] T368;
  wire[31:0] T340;
  wire T341;
  wire T342;
  wire T343;
  wire[31:0] T369;
  wire T370;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  reg  valid;
  wire dcmp_io_a_eq_b;
  wire dcmp_io_a_lt_b;
  wire dcmp_io_a_eq_b_invalid;
  wire dcmp_io_a_lt_b_invalid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_rm = {1{$random}};
    in_cmd = {1{$random}};
    in_typ = {1{$random}};
    in_single = {1{$random}};
    valid = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T22 ? T2 : T1;
  assign T1 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T2 = {T21, T3};
  assign T3 = {T10, T4};
  assign T4 = T7 | T5;
  assign T5 = T6 << 5'h1d;
  assign T6 = io_in_bits_in2[5'h16:1'h0];
  assign T7 = 52'h0 - T352;
  assign T352 = {51'h0, T8};
  assign T8 = T9 == 3'h7;
  assign T9 = io_in_bits_in2[5'h1f:5'h1d];
  assign T10 = T20 ? T354 : T11;
  assign T11 = T18 ? T353 : T12;
  assign T12 = T16 ? T15 : T13;
  assign T13 = T14 ? 12'hc00 : 12'he00;
  assign T14 = T9 < 3'h7;
  assign T15 = {4'h8, T19};
  assign T19 = io_in_bits_in2[5'h1e:5'h17];
  assign T16 = T9 < 3'h6;
  assign T353 = {1'h0, T17};
  assign T17 = {3'h7, T19};
  assign T18 = T9 < 3'h4;
  assign T354 = {4'h0, T19};
  assign T20 = T9 < 3'h1;
  assign T21 = io_in_bits_in2[6'h20:6'h20];
  assign T22 = io_in_valid & T23;
  assign T23 = T27 & T24;
  assign T24 = T25 == 1'h0;
  assign T25 = T26 == 5'hc;
  assign T26 = io_in_bits_cmd & 5'hc;
  assign T27 = io_in_bits_single & T28;
  assign T28 = io_in_bits_ldst ^ 1'h1;
  assign T29 = T22 ? T31 : T30;
  assign T30 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T31 = {T50, T32};
  assign T32 = {T39, T33};
  assign T33 = T36 | T34;
  assign T34 = T35 << 5'h1d;
  assign T35 = io_in_bits_in1[5'h16:1'h0];
  assign T36 = 52'h0 - T355;
  assign T355 = {51'h0, T37};
  assign T37 = T38 == 3'h7;
  assign T38 = io_in_bits_in1[5'h1f:5'h1d];
  assign T39 = T49 ? T357 : T40;
  assign T40 = T47 ? T356 : T41;
  assign T41 = T45 ? T44 : T42;
  assign T42 = T43 ? 12'hc00 : 12'he00;
  assign T43 = T38 < 3'h7;
  assign T44 = {4'h8, T48};
  assign T48 = io_in_bits_in1[5'h1e:5'h17];
  assign T45 = T38 < 3'h6;
  assign T356 = {1'h0, T46};
  assign T46 = {3'h7, T48};
  assign T47 = T38 < 3'h4;
  assign T357 = {4'h0, T48};
  assign T49 = T38 < 3'h1;
  assign T50 = io_in_bits_in1[6'h20:6'h20];
  assign io_out_bits_exc = T51;
  assign T51 = T150 ? T61 : T52;
  assign T52 = T58 ? dcmp_exc : 5'h0;
  assign dcmp_exc = T53 << 3'h4;
  assign T53 = T54 != 3'h0;
  assign T54 = T56 & T358;
  assign T358 = {1'h0, T55};
  assign T55 = {dcmp_io_a_lt_b_invalid, dcmp_io_a_eq_b_invalid};
  assign T56 = ~ in_rm;
  assign T57 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T58 = T59 == 5'h4;
  assign T59 = in_cmd & 5'hc;
  assign T60 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T61 = {T80, T62};
  assign T62 = {3'h0, T63};
  assign T63 = T65 & T64;
  assign T64 = T80 ^ 1'h1;
  assign T65 = T66 != 2'h0;
  assign T66 = T67[1'h1:1'h0];
  assign T67 = {T79, T68};
  assign T68 = T69 != 51'h0;
  assign T69 = T70[6'h32:1'h0];
  assign T70 = T76 << T71;
  assign T71 = T74 ? 6'h0 : T72;
  assign T72 = T73[3'h5:1'h0];
  assign T73 = in_in1[6'h3f:6'h34];
  assign T74 = T75 ^ 1'h1;
  assign T75 = T73[4'hb:4'hb];
  assign T76 = {T78, T77};
  assign T77 = in_in1[6'h33:1'h0];
  assign T78 = T74 ^ 1'h1;
  assign T79 = T70[6'h34:6'h33];
  assign T80 = T148 | T81;
  assign T81 = T147 ? T141 : T82;
  assign T82 = T140 ? T134 : T83;
  assign T83 = T131 ? T125 : T84;
  assign T84 = T74 ? 1'h0 : T85;
  assign T85 = T124 ? T120 : T86;
  assign T86 = T119 ? T89 : T87;
  assign T87 = 11'h40 <= T88;
  assign T88 = T73[4'ha:1'h0];
  assign T89 = T92 | T90;
  assign T90 = T91 != 64'h0;
  assign T91 = T70[7'h73:6'h34];
  assign T92 = T118 | T93;
  assign T93 = T117 ? T106 : T94;
  assign T94 = T105 ? T104 : T95;
  assign T95 = T103 ? T96 : 1'h0;
  assign T96 = T101 & T97;
  assign T97 = T74 ? T98 : T65;
  assign T98 = T99 ^ 1'h1;
  assign T99 = T100 == 3'h0;
  assign T100 = T73[4'hb:4'h9];
  assign T101 = T102 ^ 1'h1;
  assign T102 = in_in1[7'h40:7'h40];
  assign T103 = in_rm == 3'h3;
  assign T104 = T102 & T97;
  assign T105 = in_rm == 3'h2;
  assign T106 = T74 ? T112 : T107;
  assign T107 = T110 | T108;
  assign T108 = T109 == 2'h3;
  assign T109 = T67[1'h1:1'h0];
  assign T110 = T111 == 2'h3;
  assign T111 = T67[2'h2:1'h1];
  assign T112 = T113 & T65;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T116 == 11'h7ff;
  assign T116 = T73[4'ha:1'h0];
  assign T117 = in_rm == 3'h0;
  assign T118 = T102 ^ 1'h1;
  assign T119 = T88 == 11'h3f;
  assign T120 = T123 & T121;
  assign T121 = T93 & T122;
  assign T122 = T91 == 64'hffffffffffffffff;
  assign T123 = T102 ^ 1'h1;
  assign T124 = T88 == 11'h3e;
  assign T125 = T74 ? T130 : T126;
  assign T126 = T102 | T127;
  assign T127 = T129 ? T121 : T128;
  assign T128 = 11'h40 <= T88;
  assign T129 = T88 == 11'h3f;
  assign T130 = T102 & T93;
  assign T131 = T132 == 2'h2;
  assign T132 = in_typ ^ 2'h1;
  assign T133 = io_in_valid ? io_in_bits_typ : in_typ;
  assign T134 = T74 ? 1'h0 : T135;
  assign T135 = T139 ? T120 : T136;
  assign T136 = T138 ? T89 : T137;
  assign T137 = 11'h20 <= T88;
  assign T138 = T88 == 11'h1f;
  assign T139 = T88 == 11'h1e;
  assign T140 = T132 == 2'h1;
  assign T141 = T74 ? T146 : T142;
  assign T142 = T102 | T143;
  assign T143 = T145 ? T121 : T144;
  assign T144 = 11'h20 <= T88;
  assign T145 = T88 == 11'h1f;
  assign T146 = T102 & T93;
  assign T147 = T132 == 2'h0;
  assign T148 = T149 == 2'h3;
  assign T149 = T73[4'hb:4'ha];
  assign T150 = T151 == 5'h8;
  assign T151 = in_cmd & 5'hc;
  assign io_out_bits_toint = T152;
  assign T152 = T150 ? T327 : T153;
  assign T153 = T58 ? T363 : T154;
  assign T154 = T323 ? T362 : unrec_out;
  assign unrec_out = in_single ? T190 : unrec_d;
  assign unrec_d = {T189, T155};
  assign T155 = {T185, T156};
  assign T156 = T173 ? T172 : T157;
  assign T157 = T164 ? T158 : 52'h0;
  assign T158 = T159[6'h33:1'h0];
  assign T159 = T163 >> T160;
  assign T160 = 6'h2 - T161;
  assign T161 = T162[3'h5:1'h0];
  assign T162 = in_in1[6'h3f:6'h34];
  assign T163 = {1'h1, T172};
  assign T164 = T170 | T165;
  assign T165 = T168 & T166;
  assign T166 = T167 < 10'h2;
  assign T167 = T162[4'h9:1'h0];
  assign T168 = T169 == 2'h1;
  assign T169 = T162[4'hb:4'ha];
  assign T170 = T171 == 3'h1;
  assign T171 = T162[4'hb:4'h9];
  assign T172 = in_in1[6'h33:1'h0];
  assign T173 = T178 | T174;
  assign T174 = T176 & T175;
  assign T175 = T162[4'h9:4'h9];
  assign T176 = T177 == 2'h3;
  assign T177 = T162[4'hb:4'ha];
  assign T178 = T181 | T179;
  assign T179 = T180 == 2'h2;
  assign T180 = T162[4'hb:4'ha];
  assign T181 = T183 & T182;
  assign T182 = T166 ^ 1'h1;
  assign T183 = T184 == 2'h1;
  assign T184 = T162[4'hb:4'ha];
  assign T185 = T178 ? T187 : T186;
  assign T186 = 11'h0 - T359;
  assign T359 = {10'h0, T176};
  assign T187 = T188 - 11'h401;
  assign T188 = T162[4'ha:1'h0];
  assign T189 = in_in1[7'h40:7'h40];
  assign T190 = {T226, unrec_s};
  assign unrec_s = {T225, T191};
  assign T191 = {T221, T192};
  assign T192 = T209 ? T208 : T193;
  assign T193 = T200 ? T194 : 23'h0;
  assign T194 = T195[5'h16:1'h0];
  assign T195 = T199 >> T196;
  assign T196 = 5'h2 - T197;
  assign T197 = T198[3'h4:1'h0];
  assign T198 = in_in1[5'h1f:5'h17];
  assign T199 = {1'h1, T208};
  assign T200 = T206 | T201;
  assign T201 = T204 & T202;
  assign T202 = T203 < 7'h2;
  assign T203 = T198[3'h6:1'h0];
  assign T204 = T205 == 2'h1;
  assign T205 = T198[4'h8:3'h7];
  assign T206 = T207 == 3'h1;
  assign T207 = T198[4'h8:3'h6];
  assign T208 = in_in1[5'h16:1'h0];
  assign T209 = T214 | T210;
  assign T210 = T212 & T211;
  assign T211 = T198[3'h6:3'h6];
  assign T212 = T213 == 2'h3;
  assign T213 = T198[4'h8:3'h7];
  assign T214 = T217 | T215;
  assign T215 = T216 == 2'h2;
  assign T216 = T198[4'h8:3'h7];
  assign T217 = T219 & T218;
  assign T218 = T202 ^ 1'h1;
  assign T219 = T220 == 2'h1;
  assign T220 = T198[4'h8:3'h7];
  assign T221 = T214 ? T223 : T222;
  assign T222 = 8'h0 - T360;
  assign T360 = {7'h0, T212};
  assign T223 = T224 - 8'h81;
  assign T224 = T198[3'h7:1'h0];
  assign T225 = in_in1[6'h20:6'h20];
  assign T226 = 32'h0 - T361;
  assign T361 = {31'h0, T227};
  assign T227 = unrec_s[5'h1f:5'h1f];
  assign T228 = io_in_valid ? io_in_bits_single : in_single;
  assign T362 = {54'h0, classify_out};
  assign classify_out = in_single ? classify_s : classify_d;
  assign classify_d = {T259, T229};
  assign T229 = {T254, T230};
  assign T230 = {T249, T231};
  assign T231 = {T241, T232};
  assign T232 = T234 & T233;
  assign T233 = in_in1[7'h40:7'h40];
  assign T234 = T238 & T235;
  assign T235 = T236 ^ 1'h1;
  assign T236 = T237[4'h9:4'h9];
  assign T237 = in_in1[6'h3f:6'h34];
  assign T238 = T239 == 2'h3;
  assign T239 = T240[2'h2:1'h1];
  assign T240 = T237[4'hb:4'h9];
  assign T241 = T242 & T233;
  assign T242 = T244 | T243;
  assign T243 = T239 == 2'h2;
  assign T244 = T248 & T245;
  assign T245 = T246 ^ 1'h1;
  assign T246 = T247 < 10'h2;
  assign T247 = T237[4'h9:1'h0];
  assign T248 = T239 == 2'h1;
  assign T249 = T250 & T233;
  assign T250 = T253 | T251;
  assign T251 = T252 & T246;
  assign T252 = T239 == 2'h1;
  assign T253 = T240 == 3'h1;
  assign T254 = {T257, T255};
  assign T255 = T256 & T233;
  assign T256 = T240 == 3'h0;
  assign T257 = T256 & T258;
  assign T258 = T233 ^ 1'h1;
  assign T259 = {T268, T260};
  assign T260 = {T266, T261};
  assign T261 = {T264, T262};
  assign T262 = T250 & T263;
  assign T263 = T233 ^ 1'h1;
  assign T264 = T242 & T265;
  assign T265 = T233 ^ 1'h1;
  assign T266 = T234 & T267;
  assign T267 = T233 ^ 1'h1;
  assign T268 = {T274, T269};
  assign T269 = T273 & T270;
  assign T270 = T271 ^ 1'h1;
  assign T271 = T272[6'h33:6'h33];
  assign T272 = in_in1[6'h33:1'h0];
  assign T273 = T240 == 3'h7;
  assign T274 = T273 & T275;
  assign T275 = T272[6'h33:6'h33];
  assign classify_s = {T306, T276};
  assign T276 = {T301, T277};
  assign T277 = {T296, T278};
  assign T278 = {T288, T279};
  assign T279 = T281 & T280;
  assign T280 = in_in1[6'h20:6'h20];
  assign T281 = T285 & T282;
  assign T282 = T283 ^ 1'h1;
  assign T283 = T284[3'h6:3'h6];
  assign T284 = in_in1[5'h1f:5'h17];
  assign T285 = T286 == 2'h3;
  assign T286 = T287[2'h2:1'h1];
  assign T287 = T284[4'h8:3'h6];
  assign T288 = T289 & T280;
  assign T289 = T291 | T290;
  assign T290 = T286 == 2'h2;
  assign T291 = T295 & T292;
  assign T292 = T293 ^ 1'h1;
  assign T293 = T294 < 7'h2;
  assign T294 = T284[3'h6:1'h0];
  assign T295 = T286 == 2'h1;
  assign T296 = T297 & T280;
  assign T297 = T300 | T298;
  assign T298 = T299 & T293;
  assign T299 = T286 == 2'h1;
  assign T300 = T287 == 3'h1;
  assign T301 = {T304, T302};
  assign T302 = T303 & T280;
  assign T303 = T287 == 3'h0;
  assign T304 = T303 & T305;
  assign T305 = T280 ^ 1'h1;
  assign T306 = {T315, T307};
  assign T307 = {T313, T308};
  assign T308 = {T311, T309};
  assign T309 = T297 & T310;
  assign T310 = T280 ^ 1'h1;
  assign T311 = T289 & T312;
  assign T312 = T280 ^ 1'h1;
  assign T313 = T281 & T314;
  assign T314 = T280 ^ 1'h1;
  assign T315 = {T321, T316};
  assign T316 = T320 & T317;
  assign T317 = T318 ^ 1'h1;
  assign T318 = T319[5'h16:5'h16];
  assign T319 = in_in1[5'h16:1'h0];
  assign T320 = T287 == 3'h7;
  assign T321 = T320 & T322;
  assign T322 = T319[5'h16:5'h16];
  assign T323 = in_rm[1'h0:1'h0];
  assign T363 = {63'h0, dcmp_out};
  assign dcmp_out = T324 != 3'h0;
  assign T324 = T326 & T364;
  assign T364 = {1'h0, T325};
  assign T325 = {dcmp_io_a_lt_b, dcmp_io_a_eq_b};
  assign T326 = ~ in_rm;
  assign T327 = T351 ? T330 : T365;
  assign T365 = {T366, T328};
  assign T328 = T329;
  assign T329 = T330[5'h1f:1'h0];
  assign T366 = T367 ? 32'hffffffff : 32'h0;
  assign T367 = T328[5'h1f:5'h1f];
  assign T330 = T80 ? T337 : T331;
  assign T331 = T332;
  assign T332 = T336 ? T335 : T333;
  assign T333 = T102 ? T334 : T91;
  assign T334 = ~ T91;
  assign T335 = T333 + 64'h1;
  assign T336 = T93 ^ T102;
  assign T337 = T349 ? 64'h8000000000000000 : T338;
  assign T338 = T347 ? 64'hffffffff80000000 : T339;
  assign T339 = T344 ? 64'h7fffffffffffffff : T368;
  assign T368 = {T369, T340};
  assign T340 = T341 ? 32'h7fffffff : 32'hffffffff;
  assign T341 = T343 & T342;
  assign T342 = T102 ^ 1'h1;
  assign T343 = T132 == 2'h1;
  assign T369 = T370 ? 32'hffffffff : 32'h0;
  assign T370 = T340[5'h1f:5'h1f];
  assign T344 = T346 & T345;
  assign T345 = T102 ^ 1'h1;
  assign T346 = T132 == 2'h3;
  assign T347 = T348 & T102;
  assign T348 = T132 == 2'h1;
  assign T349 = T350 & T102;
  assign T350 = T132 == 2'h3;
  assign T351 = in_typ[1'h1:1'h1];
  assign io_out_bits_store = unrec_out;
  assign io_out_bits_lt = dcmp_io_a_lt_b;
  assign io_out_valid = valid;
  recodedFloatNCompare dcmp(
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_a_eq_b( dcmp_io_a_eq_b ),
       .io_a_lt_b( dcmp_io_a_lt_b ),
       .io_a_eq_b_invalid( dcmp_io_a_eq_b_invalid ),
       .io_a_lt_b_invalid( dcmp_io_a_lt_b_invalid )
  );

  always @(posedge clk) begin
    if(T22) begin
      in_in2 <= T2;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(T22) begin
      in_in1 <= T31;
    end else if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      in_single <= io_in_bits_single;
    end
    valid <= io_in_valid;
  end
endmodule

module IntToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  reg [4:0] R0;
  wire[4:0] T1;
  reg [4:0] R2;
  wire[4:0] T3;
  wire[4:0] mux_exc;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[1:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[38:0] T12;
  wire[126:0] T13;
  wire[5:0] T14;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[5:0] T210;
  wire[5:0] T211;
  wire[5:0] T212;
  wire[5:0] T213;
  wire[5:0] T214;
  wire[5:0] T215;
  wire[5:0] T216;
  wire[5:0] T217;
  wire[5:0] T218;
  wire[5:0] T219;
  wire[5:0] T220;
  wire[5:0] T221;
  wire[5:0] T222;
  wire[5:0] T223;
  wire[5:0] T224;
  wire[5:0] T225;
  wire[5:0] T226;
  wire[5:0] T227;
  wire[5:0] T228;
  wire[5:0] T229;
  wire[5:0] T230;
  wire[5:0] T231;
  wire[5:0] T232;
  wire[5:0] T233;
  wire[5:0] T234;
  wire[5:0] T235;
  wire[5:0] T236;
  wire[5:0] T237;
  wire[5:0] T238;
  wire[4:0] T239;
  wire[4:0] T240;
  wire[4:0] T241;
  wire[4:0] T242;
  wire[4:0] T243;
  wire[4:0] T244;
  wire[4:0] T245;
  wire[4:0] T246;
  wire[4:0] T247;
  wire[4:0] T248;
  wire[4:0] T249;
  wire[4:0] T250;
  wire[4:0] T251;
  wire[4:0] T252;
  wire[4:0] T253;
  wire[4:0] T254;
  wire[3:0] T255;
  wire[3:0] T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[3:0] T262;
  wire[2:0] T263;
  wire[2:0] T264;
  wire[2:0] T265;
  wire[2:0] T266;
  wire[1:0] T267;
  wire[1:0] T268;
  wire T269;
  wire[63:0] T16;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[63:0] T17;
  wire[63:0] T332;
  wire[31:0] T18;
  wire[63:0] T19;
  wire[63:0] T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire[63:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  reg [1:0] R29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  reg  R38;
  wire T39;
  wire T40;
  wire[4:0] T41;
  reg [4:0] R42;
  wire[4:0] T43;
  wire[4:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire[2:0] T48;
  wire T49;
  wire[9:0] T50;
  wire[126:0] T51;
  wire[5:0] T52;
  wire[5:0] T333;
  wire[5:0] T334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[5:0] T338;
  wire[5:0] T339;
  wire[5:0] T340;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[5:0] T343;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[5:0] T349;
  wire[5:0] T350;
  wire[5:0] T351;
  wire[5:0] T352;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[5:0] T357;
  wire[5:0] T358;
  wire[5:0] T359;
  wire[5:0] T360;
  wire[5:0] T361;
  wire[5:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[4:0] T365;
  wire[4:0] T366;
  wire[4:0] T367;
  wire[4:0] T368;
  wire[4:0] T369;
  wire[4:0] T370;
  wire[4:0] T371;
  wire[4:0] T372;
  wire[4:0] T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire[4:0] T377;
  wire[4:0] T378;
  wire[4:0] T379;
  wire[4:0] T380;
  wire[3:0] T381;
  wire[3:0] T382;
  wire[3:0] T383;
  wire[3:0] T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[2:0] T389;
  wire[2:0] T390;
  wire[2:0] T391;
  wire[2:0] T392;
  wire[1:0] T393;
  wire[1:0] T394;
  wire T395;
  wire[63:0] T54;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire[63:0] T55;
  wire[63:0] T458;
  wire[31:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[1:0] T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T459;
  reg  R74;
  wire T460;
  reg [64:0] R75;
  wire[64:0] T76;
  reg [64:0] R77;
  wire[64:0] T78;
  wire[64:0] mux_data;
  wire[64:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[64:0] T82;
  wire[63:0] T83;
  wire[51:0] T84;
  wire[51:0] T85;
  wire[51:0] T86;
  wire[126:0] T87;
  wire[5:0] T88;
  wire[5:0] T461;
  wire[5:0] T462;
  wire[5:0] T463;
  wire[5:0] T464;
  wire[5:0] T465;
  wire[5:0] T466;
  wire[5:0] T467;
  wire[5:0] T468;
  wire[5:0] T469;
  wire[5:0] T470;
  wire[5:0] T471;
  wire[5:0] T472;
  wire[5:0] T473;
  wire[5:0] T474;
  wire[5:0] T475;
  wire[5:0] T476;
  wire[5:0] T477;
  wire[5:0] T478;
  wire[5:0] T479;
  wire[5:0] T480;
  wire[5:0] T481;
  wire[5:0] T482;
  wire[5:0] T483;
  wire[5:0] T484;
  wire[5:0] T485;
  wire[5:0] T486;
  wire[5:0] T487;
  wire[5:0] T488;
  wire[5:0] T489;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[5:0] T492;
  wire[4:0] T493;
  wire[4:0] T494;
  wire[4:0] T495;
  wire[4:0] T496;
  wire[4:0] T497;
  wire[4:0] T498;
  wire[4:0] T499;
  wire[4:0] T500;
  wire[4:0] T501;
  wire[4:0] T502;
  wire[4:0] T503;
  wire[4:0] T504;
  wire[4:0] T505;
  wire[4:0] T506;
  wire[4:0] T507;
  wire[4:0] T508;
  wire[3:0] T509;
  wire[3:0] T510;
  wire[3:0] T511;
  wire[3:0] T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[3:0] T516;
  wire[2:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire[2:0] T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire T523;
  wire[63:0] T90;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[63:0] T91;
  wire T92;
  wire[10:0] T93;
  wire[11:0] T94;
  wire[11:0] T586;
  wire[9:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[11:0] T101;
  wire[11:0] T587;
  wire[10:0] T102;
  wire[10:0] T103;
  wire[10:0] T588;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[11:0] T108;
  wire[11:0] T589;
  wire[11:0] T109;
  wire[11:0] T110;
  wire[5:0] T111;
  wire T112;
  wire[64:0] T113;
  wire[32:0] T114;
  wire[31:0] T115;
  wire[22:0] T116;
  wire[22:0] T117;
  wire[22:0] T118;
  wire[62:0] T119;
  wire[4:0] T120;
  wire[4:0] T590;
  wire[4:0] T591;
  wire[4:0] T592;
  wire[4:0] T593;
  wire[4:0] T594;
  wire[4:0] T595;
  wire[4:0] T596;
  wire[4:0] T597;
  wire[4:0] T598;
  wire[4:0] T599;
  wire[4:0] T600;
  wire[4:0] T601;
  wire[4:0] T602;
  wire[4:0] T603;
  wire[4:0] T604;
  wire[4:0] T605;
  wire[3:0] T606;
  wire[3:0] T607;
  wire[3:0] T608;
  wire[3:0] T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[3:0] T612;
  wire[3:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire[2:0] T616;
  wire[2:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire T620;
  wire[31:0] T122;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire[31:0] T123;
  wire T124;
  wire[7:0] T125;
  wire[8:0] T126;
  wire[8:0] T651;
  wire[6:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  wire[8:0] T133;
  wire[8:0] T652;
  wire[7:0] T134;
  wire[7:0] T135;
  wire[7:0] T653;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire[8:0] T140;
  wire[8:0] T654;
  wire[8:0] T141;
  wire[8:0] T142;
  wire[4:0] T143;
  wire T144;
  wire[64:0] T145;
  wire[32:0] T146;
  wire[31:0] T147;
  wire[22:0] T148;
  wire[24:0] T149;
  wire[24:0] T150;
  wire[23:0] T151;
  wire[24:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  reg [2:0] R159;
  wire[2:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire[1:0] T167;
  wire T168;
  wire[8:0] T169;
  wire[7:0] T170;
  wire[7:0] T171;
  wire[7:0] T655;
  wire T172;
  wire[7:0] T173;
  wire[6:0] T174;
  wire[5:0] T175;
  wire T176;
  wire[64:0] T177;
  wire[63:0] T178;
  wire[51:0] T179;
  wire[53:0] T180;
  wire[53:0] T181;
  wire[52:0] T182;
  wire[53:0] T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[1:0] T194;
  wire T195;
  wire[1:0] T196;
  wire T197;
  wire[11:0] T198;
  wire[10:0] T199;
  wire[10:0] T200;
  wire[10:0] T656;
  wire T201;
  wire[10:0] T202;
  wire[9:0] T203;
  wire[5:0] T204;
  wire T205;
  reg  R206;
  wire T657;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R2 = {1{$random}};
    R21 = {3{$random}};
    R29 = {1{$random}};
    R38 = {1{$random}};
    R42 = {1{$random}};
    R73 = {1{$random}};
    R74 = {1{$random}};
    R75 = {3{$random}};
    R77 = {3{$random}};
    R159 = {1{$random}};
    R206 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R74 ? R2 : R0;
  assign T3 = R73 ? mux_exc : R2;
  assign mux_exc = T4;
  assign T4 = T71 ? T44 : T5;
  assign T5 = T37 ? T6 : 5'h0;
  assign T6 = {3'h0, T7};
  assign T7 = {1'h0, T8};
  assign T8 = T9 != 2'h0;
  assign T9 = T10[1'h1:1'h0];
  assign T10 = {T36, T11};
  assign T11 = T12 != 39'h0;
  assign T12 = T13[6'h26:1'h0];
  assign T13 = T17 << T14;
  assign T14 = ~ T207;
  assign T207 = T331 ? 6'h3f : T208;
  assign T208 = T330 ? 6'h3e : T209;
  assign T209 = T329 ? 6'h3d : T210;
  assign T210 = T328 ? 6'h3c : T211;
  assign T211 = T327 ? 6'h3b : T212;
  assign T212 = T326 ? 6'h3a : T213;
  assign T213 = T325 ? 6'h39 : T214;
  assign T214 = T324 ? 6'h38 : T215;
  assign T215 = T323 ? 6'h37 : T216;
  assign T216 = T322 ? 6'h36 : T217;
  assign T217 = T321 ? 6'h35 : T218;
  assign T218 = T320 ? 6'h34 : T219;
  assign T219 = T319 ? 6'h33 : T220;
  assign T220 = T318 ? 6'h32 : T221;
  assign T221 = T317 ? 6'h31 : T222;
  assign T222 = T316 ? 6'h30 : T223;
  assign T223 = T315 ? 6'h2f : T224;
  assign T224 = T314 ? 6'h2e : T225;
  assign T225 = T313 ? 6'h2d : T226;
  assign T226 = T312 ? 6'h2c : T227;
  assign T227 = T311 ? 6'h2b : T228;
  assign T228 = T310 ? 6'h2a : T229;
  assign T229 = T309 ? 6'h29 : T230;
  assign T230 = T308 ? 6'h28 : T231;
  assign T231 = T307 ? 6'h27 : T232;
  assign T232 = T306 ? 6'h26 : T233;
  assign T233 = T305 ? 6'h25 : T234;
  assign T234 = T304 ? 6'h24 : T235;
  assign T235 = T303 ? 6'h23 : T236;
  assign T236 = T302 ? 6'h22 : T237;
  assign T237 = T301 ? 6'h21 : T238;
  assign T238 = T300 ? 6'h20 : T239;
  assign T239 = T299 ? 5'h1f : T240;
  assign T240 = T298 ? 5'h1e : T241;
  assign T241 = T297 ? 5'h1d : T242;
  assign T242 = T296 ? 5'h1c : T243;
  assign T243 = T295 ? 5'h1b : T244;
  assign T244 = T294 ? 5'h1a : T245;
  assign T245 = T293 ? 5'h19 : T246;
  assign T246 = T292 ? 5'h18 : T247;
  assign T247 = T291 ? 5'h17 : T248;
  assign T248 = T290 ? 5'h16 : T249;
  assign T249 = T289 ? 5'h15 : T250;
  assign T250 = T288 ? 5'h14 : T251;
  assign T251 = T287 ? 5'h13 : T252;
  assign T252 = T286 ? 5'h12 : T253;
  assign T253 = T285 ? 5'h11 : T254;
  assign T254 = T284 ? 5'h10 : T255;
  assign T255 = T283 ? 4'hf : T256;
  assign T256 = T282 ? 4'he : T257;
  assign T257 = T281 ? 4'hd : T258;
  assign T258 = T280 ? 4'hc : T259;
  assign T259 = T279 ? 4'hb : T260;
  assign T260 = T278 ? 4'ha : T261;
  assign T261 = T277 ? 4'h9 : T262;
  assign T262 = T276 ? 4'h8 : T263;
  assign T263 = T275 ? 3'h7 : T264;
  assign T264 = T274 ? 3'h6 : T265;
  assign T265 = T273 ? 3'h5 : T266;
  assign T266 = T272 ? 3'h4 : T267;
  assign T267 = T271 ? 2'h3 : T268;
  assign T268 = T270 ? 2'h2 : T269;
  assign T269 = T16[1'h1:1'h1];
  assign T16 = T17[6'h3f:1'h0];
  assign T270 = T16[2'h2:2'h2];
  assign T271 = T16[2'h3:2'h3];
  assign T272 = T16[3'h4:3'h4];
  assign T273 = T16[3'h5:3'h5];
  assign T274 = T16[3'h6:3'h6];
  assign T275 = T16[3'h7:3'h7];
  assign T276 = T16[4'h8:4'h8];
  assign T277 = T16[4'h9:4'h9];
  assign T278 = T16[4'ha:4'ha];
  assign T279 = T16[4'hb:4'hb];
  assign T280 = T16[4'hc:4'hc];
  assign T281 = T16[4'hd:4'hd];
  assign T282 = T16[4'he:4'he];
  assign T283 = T16[4'hf:4'hf];
  assign T284 = T16[5'h10:5'h10];
  assign T285 = T16[5'h11:5'h11];
  assign T286 = T16[5'h12:5'h12];
  assign T287 = T16[5'h13:5'h13];
  assign T288 = T16[5'h14:5'h14];
  assign T289 = T16[5'h15:5'h15];
  assign T290 = T16[5'h16:5'h16];
  assign T291 = T16[5'h17:5'h17];
  assign T292 = T16[5'h18:5'h18];
  assign T293 = T16[5'h19:5'h19];
  assign T294 = T16[5'h1a:5'h1a];
  assign T295 = T16[5'h1b:5'h1b];
  assign T296 = T16[5'h1c:5'h1c];
  assign T297 = T16[5'h1d:5'h1d];
  assign T298 = T16[5'h1e:5'h1e];
  assign T299 = T16[5'h1f:5'h1f];
  assign T300 = T16[6'h20:6'h20];
  assign T301 = T16[6'h21:6'h21];
  assign T302 = T16[6'h22:6'h22];
  assign T303 = T16[6'h23:6'h23];
  assign T304 = T16[6'h24:6'h24];
  assign T305 = T16[6'h25:6'h25];
  assign T306 = T16[6'h26:6'h26];
  assign T307 = T16[6'h27:6'h27];
  assign T308 = T16[6'h28:6'h28];
  assign T309 = T16[6'h29:6'h29];
  assign T310 = T16[6'h2a:6'h2a];
  assign T311 = T16[6'h2b:6'h2b];
  assign T312 = T16[6'h2c:6'h2c];
  assign T313 = T16[6'h2d:6'h2d];
  assign T314 = T16[6'h2e:6'h2e];
  assign T315 = T16[6'h2f:6'h2f];
  assign T316 = T16[6'h30:6'h30];
  assign T317 = T16[6'h31:6'h31];
  assign T318 = T16[6'h32:6'h32];
  assign T319 = T16[6'h33:6'h33];
  assign T320 = T16[6'h34:6'h34];
  assign T321 = T16[6'h35:6'h35];
  assign T322 = T16[6'h36:6'h36];
  assign T323 = T16[6'h37:6'h37];
  assign T324 = T16[6'h38:6'h38];
  assign T325 = T16[6'h39:6'h39];
  assign T326 = T16[6'h3a:6'h3a];
  assign T327 = T16[6'h3b:6'h3b];
  assign T328 = T16[6'h3c:6'h3c];
  assign T329 = T16[6'h3d:6'h3d];
  assign T330 = T16[6'h3e:6'h3e];
  assign T331 = T16[6'h3f:6'h3f];
  assign T17 = T33 ? T19 : T332;
  assign T332 = {32'h0, T18};
  assign T18 = T19[5'h1f:1'h0];
  assign T19 = T24 ? T23 : T20;
  assign T20 = R21[6'h3f:1'h0];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = 64'h0 - T20;
  assign T24 = T32 ? T31 : T25;
  assign T25 = T27 ? T26 : 1'h0;
  assign T26 = T20[6'h3f:6'h3f];
  assign T27 = T28 == 2'h3;
  assign T28 = R29 ^ 2'h1;
  assign T30 = io_in_valid ? io_in_bits_typ : R29;
  assign T31 = T20[5'h1f:5'h1f];
  assign T32 = T28 == 2'h1;
  assign T33 = T35 | T34;
  assign T34 = T28 == 2'h2;
  assign T35 = T28 == 2'h3;
  assign T36 = T13[6'h28:6'h27];
  assign T37 = T40 & R38;
  assign T39 = io_in_valid ? io_in_bits_single : R38;
  assign T40 = T41 == 5'h0;
  assign T41 = R42 & 5'h4;
  assign T43 = io_in_valid ? io_in_bits_cmd : R42;
  assign T44 = {3'h0, T45};
  assign T45 = {1'h0, T46};
  assign T46 = T47 != 2'h0;
  assign T47 = T48[1'h1:1'h0];
  assign T48 = {T70, T49};
  assign T49 = T50 != 10'h0;
  assign T50 = T51[4'h9:1'h0];
  assign T51 = T55 << T52;
  assign T52 = ~ T333;
  assign T333 = T457 ? 6'h3f : T334;
  assign T334 = T456 ? 6'h3e : T335;
  assign T335 = T455 ? 6'h3d : T336;
  assign T336 = T454 ? 6'h3c : T337;
  assign T337 = T453 ? 6'h3b : T338;
  assign T338 = T452 ? 6'h3a : T339;
  assign T339 = T451 ? 6'h39 : T340;
  assign T340 = T450 ? 6'h38 : T341;
  assign T341 = T449 ? 6'h37 : T342;
  assign T342 = T448 ? 6'h36 : T343;
  assign T343 = T447 ? 6'h35 : T344;
  assign T344 = T446 ? 6'h34 : T345;
  assign T345 = T445 ? 6'h33 : T346;
  assign T346 = T444 ? 6'h32 : T347;
  assign T347 = T443 ? 6'h31 : T348;
  assign T348 = T442 ? 6'h30 : T349;
  assign T349 = T441 ? 6'h2f : T350;
  assign T350 = T440 ? 6'h2e : T351;
  assign T351 = T439 ? 6'h2d : T352;
  assign T352 = T438 ? 6'h2c : T353;
  assign T353 = T437 ? 6'h2b : T354;
  assign T354 = T436 ? 6'h2a : T355;
  assign T355 = T435 ? 6'h29 : T356;
  assign T356 = T434 ? 6'h28 : T357;
  assign T357 = T433 ? 6'h27 : T358;
  assign T358 = T432 ? 6'h26 : T359;
  assign T359 = T431 ? 6'h25 : T360;
  assign T360 = T430 ? 6'h24 : T361;
  assign T361 = T429 ? 6'h23 : T362;
  assign T362 = T428 ? 6'h22 : T363;
  assign T363 = T427 ? 6'h21 : T364;
  assign T364 = T426 ? 6'h20 : T365;
  assign T365 = T425 ? 5'h1f : T366;
  assign T366 = T424 ? 5'h1e : T367;
  assign T367 = T423 ? 5'h1d : T368;
  assign T368 = T422 ? 5'h1c : T369;
  assign T369 = T421 ? 5'h1b : T370;
  assign T370 = T420 ? 5'h1a : T371;
  assign T371 = T419 ? 5'h19 : T372;
  assign T372 = T418 ? 5'h18 : T373;
  assign T373 = T417 ? 5'h17 : T374;
  assign T374 = T416 ? 5'h16 : T375;
  assign T375 = T415 ? 5'h15 : T376;
  assign T376 = T414 ? 5'h14 : T377;
  assign T377 = T413 ? 5'h13 : T378;
  assign T378 = T412 ? 5'h12 : T379;
  assign T379 = T411 ? 5'h11 : T380;
  assign T380 = T410 ? 5'h10 : T381;
  assign T381 = T409 ? 4'hf : T382;
  assign T382 = T408 ? 4'he : T383;
  assign T383 = T407 ? 4'hd : T384;
  assign T384 = T406 ? 4'hc : T385;
  assign T385 = T405 ? 4'hb : T386;
  assign T386 = T404 ? 4'ha : T387;
  assign T387 = T403 ? 4'h9 : T388;
  assign T388 = T402 ? 4'h8 : T389;
  assign T389 = T401 ? 3'h7 : T390;
  assign T390 = T400 ? 3'h6 : T391;
  assign T391 = T399 ? 3'h5 : T392;
  assign T392 = T398 ? 3'h4 : T393;
  assign T393 = T397 ? 2'h3 : T394;
  assign T394 = T396 ? 2'h2 : T395;
  assign T395 = T54[1'h1:1'h1];
  assign T54 = T55[6'h3f:1'h0];
  assign T396 = T54[2'h2:2'h2];
  assign T397 = T54[2'h3:2'h3];
  assign T398 = T54[3'h4:3'h4];
  assign T399 = T54[3'h5:3'h5];
  assign T400 = T54[3'h6:3'h6];
  assign T401 = T54[3'h7:3'h7];
  assign T402 = T54[4'h8:4'h8];
  assign T403 = T54[4'h9:4'h9];
  assign T404 = T54[4'ha:4'ha];
  assign T405 = T54[4'hb:4'hb];
  assign T406 = T54[4'hc:4'hc];
  assign T407 = T54[4'hd:4'hd];
  assign T408 = T54[4'he:4'he];
  assign T409 = T54[4'hf:4'hf];
  assign T410 = T54[5'h10:5'h10];
  assign T411 = T54[5'h11:5'h11];
  assign T412 = T54[5'h12:5'h12];
  assign T413 = T54[5'h13:5'h13];
  assign T414 = T54[5'h14:5'h14];
  assign T415 = T54[5'h15:5'h15];
  assign T416 = T54[5'h16:5'h16];
  assign T417 = T54[5'h17:5'h17];
  assign T418 = T54[5'h18:5'h18];
  assign T419 = T54[5'h19:5'h19];
  assign T420 = T54[5'h1a:5'h1a];
  assign T421 = T54[5'h1b:5'h1b];
  assign T422 = T54[5'h1c:5'h1c];
  assign T423 = T54[5'h1d:5'h1d];
  assign T424 = T54[5'h1e:5'h1e];
  assign T425 = T54[5'h1f:5'h1f];
  assign T426 = T54[6'h20:6'h20];
  assign T427 = T54[6'h21:6'h21];
  assign T428 = T54[6'h22:6'h22];
  assign T429 = T54[6'h23:6'h23];
  assign T430 = T54[6'h24:6'h24];
  assign T431 = T54[6'h25:6'h25];
  assign T432 = T54[6'h26:6'h26];
  assign T433 = T54[6'h27:6'h27];
  assign T434 = T54[6'h28:6'h28];
  assign T435 = T54[6'h29:6'h29];
  assign T436 = T54[6'h2a:6'h2a];
  assign T437 = T54[6'h2b:6'h2b];
  assign T438 = T54[6'h2c:6'h2c];
  assign T439 = T54[6'h2d:6'h2d];
  assign T440 = T54[6'h2e:6'h2e];
  assign T441 = T54[6'h2f:6'h2f];
  assign T442 = T54[6'h30:6'h30];
  assign T443 = T54[6'h31:6'h31];
  assign T444 = T54[6'h32:6'h32];
  assign T445 = T54[6'h33:6'h33];
  assign T446 = T54[6'h34:6'h34];
  assign T447 = T54[6'h35:6'h35];
  assign T448 = T54[6'h36:6'h36];
  assign T449 = T54[6'h37:6'h37];
  assign T450 = T54[6'h38:6'h38];
  assign T451 = T54[6'h39:6'h39];
  assign T452 = T54[6'h3a:6'h3a];
  assign T453 = T54[6'h3b:6'h3b];
  assign T454 = T54[6'h3c:6'h3c];
  assign T455 = T54[6'h3d:6'h3d];
  assign T456 = T54[6'h3e:6'h3e];
  assign T457 = T54[6'h3f:6'h3f];
  assign T55 = T67 ? T57 : T458;
  assign T458 = {32'h0, T56};
  assign T56 = T57[5'h1f:1'h0];
  assign T57 = T60 ? T59 : T58;
  assign T58 = R21[6'h3f:1'h0];
  assign T59 = 64'h0 - T58;
  assign T60 = T66 ? T65 : T61;
  assign T61 = T63 ? T62 : 1'h0;
  assign T62 = T58[6'h3f:6'h3f];
  assign T63 = T64 == 2'h3;
  assign T64 = R29 ^ 2'h1;
  assign T65 = T58[5'h1f:5'h1f];
  assign T66 = T64 == 2'h1;
  assign T67 = T69 | T68;
  assign T68 = T64 == 2'h2;
  assign T69 = T64 == 2'h3;
  assign T70 = T51[4'hb:4'ha];
  assign T71 = T40 & T72;
  assign T72 = R38 ^ 1'h1;
  assign T459 = reset ? 1'h0 : io_in_valid;
  assign T460 = reset ? 1'h0 : R73;
  assign io_out_bits_data = R75;
  assign T76 = R74 ? R77 : R75;
  assign T78 = R73 ? mux_data : R77;
  assign mux_data = T79;
  assign T79 = T71 ? T177 : T80;
  assign T80 = T37 ? T145 : T81;
  assign T81 = R38 ? T113 : T82;
  assign T82 = {T112, T83};
  assign T83 = {T94, T84};
  assign T84 = T92 ? T86 : T85;
  assign T85 = R21[6'h33:1'h0];
  assign T86 = T87[6'h3e:4'hb];
  assign T87 = T91 << T88;
  assign T88 = ~ T461;
  assign T461 = T585 ? 6'h3f : T462;
  assign T462 = T584 ? 6'h3e : T463;
  assign T463 = T583 ? 6'h3d : T464;
  assign T464 = T582 ? 6'h3c : T465;
  assign T465 = T581 ? 6'h3b : T466;
  assign T466 = T580 ? 6'h3a : T467;
  assign T467 = T579 ? 6'h39 : T468;
  assign T468 = T578 ? 6'h38 : T469;
  assign T469 = T577 ? 6'h37 : T470;
  assign T470 = T576 ? 6'h36 : T471;
  assign T471 = T575 ? 6'h35 : T472;
  assign T472 = T574 ? 6'h34 : T473;
  assign T473 = T573 ? 6'h33 : T474;
  assign T474 = T572 ? 6'h32 : T475;
  assign T475 = T571 ? 6'h31 : T476;
  assign T476 = T570 ? 6'h30 : T477;
  assign T477 = T569 ? 6'h2f : T478;
  assign T478 = T568 ? 6'h2e : T479;
  assign T479 = T567 ? 6'h2d : T480;
  assign T480 = T566 ? 6'h2c : T481;
  assign T481 = T565 ? 6'h2b : T482;
  assign T482 = T564 ? 6'h2a : T483;
  assign T483 = T563 ? 6'h29 : T484;
  assign T484 = T562 ? 6'h28 : T485;
  assign T485 = T561 ? 6'h27 : T486;
  assign T486 = T560 ? 6'h26 : T487;
  assign T487 = T559 ? 6'h25 : T488;
  assign T488 = T558 ? 6'h24 : T489;
  assign T489 = T557 ? 6'h23 : T490;
  assign T490 = T556 ? 6'h22 : T491;
  assign T491 = T555 ? 6'h21 : T492;
  assign T492 = T554 ? 6'h20 : T493;
  assign T493 = T553 ? 5'h1f : T494;
  assign T494 = T552 ? 5'h1e : T495;
  assign T495 = T551 ? 5'h1d : T496;
  assign T496 = T550 ? 5'h1c : T497;
  assign T497 = T549 ? 5'h1b : T498;
  assign T498 = T548 ? 5'h1a : T499;
  assign T499 = T547 ? 5'h19 : T500;
  assign T500 = T546 ? 5'h18 : T501;
  assign T501 = T545 ? 5'h17 : T502;
  assign T502 = T544 ? 5'h16 : T503;
  assign T503 = T543 ? 5'h15 : T504;
  assign T504 = T542 ? 5'h14 : T505;
  assign T505 = T541 ? 5'h13 : T506;
  assign T506 = T540 ? 5'h12 : T507;
  assign T507 = T539 ? 5'h11 : T508;
  assign T508 = T538 ? 5'h10 : T509;
  assign T509 = T537 ? 4'hf : T510;
  assign T510 = T536 ? 4'he : T511;
  assign T511 = T535 ? 4'hd : T512;
  assign T512 = T534 ? 4'hc : T513;
  assign T513 = T533 ? 4'hb : T514;
  assign T514 = T532 ? 4'ha : T515;
  assign T515 = T531 ? 4'h9 : T516;
  assign T516 = T530 ? 4'h8 : T517;
  assign T517 = T529 ? 3'h7 : T518;
  assign T518 = T528 ? 3'h6 : T519;
  assign T519 = T527 ? 3'h5 : T520;
  assign T520 = T526 ? 3'h4 : T521;
  assign T521 = T525 ? 2'h3 : T522;
  assign T522 = T524 ? 2'h2 : T523;
  assign T523 = T90[1'h1:1'h1];
  assign T90 = T91[6'h3f:1'h0];
  assign T524 = T90[2'h2:2'h2];
  assign T525 = T90[2'h3:2'h3];
  assign T526 = T90[3'h4:3'h4];
  assign T527 = T90[3'h5:3'h5];
  assign T528 = T90[3'h6:3'h6];
  assign T529 = T90[3'h7:3'h7];
  assign T530 = T90[4'h8:4'h8];
  assign T531 = T90[4'h9:4'h9];
  assign T532 = T90[4'ha:4'ha];
  assign T533 = T90[4'hb:4'hb];
  assign T534 = T90[4'hc:4'hc];
  assign T535 = T90[4'hd:4'hd];
  assign T536 = T90[4'he:4'he];
  assign T537 = T90[4'hf:4'hf];
  assign T538 = T90[5'h10:5'h10];
  assign T539 = T90[5'h11:5'h11];
  assign T540 = T90[5'h12:5'h12];
  assign T541 = T90[5'h13:5'h13];
  assign T542 = T90[5'h14:5'h14];
  assign T543 = T90[5'h15:5'h15];
  assign T544 = T90[5'h16:5'h16];
  assign T545 = T90[5'h17:5'h17];
  assign T546 = T90[5'h18:5'h18];
  assign T547 = T90[5'h19:5'h19];
  assign T548 = T90[5'h1a:5'h1a];
  assign T549 = T90[5'h1b:5'h1b];
  assign T550 = T90[5'h1c:5'h1c];
  assign T551 = T90[5'h1d:5'h1d];
  assign T552 = T90[5'h1e:5'h1e];
  assign T553 = T90[5'h1f:5'h1f];
  assign T554 = T90[6'h20:6'h20];
  assign T555 = T90[6'h21:6'h21];
  assign T556 = T90[6'h22:6'h22];
  assign T557 = T90[6'h23:6'h23];
  assign T558 = T90[6'h24:6'h24];
  assign T559 = T90[6'h25:6'h25];
  assign T560 = T90[6'h26:6'h26];
  assign T561 = T90[6'h27:6'h27];
  assign T562 = T90[6'h28:6'h28];
  assign T563 = T90[6'h29:6'h29];
  assign T564 = T90[6'h2a:6'h2a];
  assign T565 = T90[6'h2b:6'h2b];
  assign T566 = T90[6'h2c:6'h2c];
  assign T567 = T90[6'h2d:6'h2d];
  assign T568 = T90[6'h2e:6'h2e];
  assign T569 = T90[6'h2f:6'h2f];
  assign T570 = T90[6'h30:6'h30];
  assign T571 = T90[6'h31:6'h31];
  assign T572 = T90[6'h32:6'h32];
  assign T573 = T90[6'h33:6'h33];
  assign T574 = T90[6'h34:6'h34];
  assign T575 = T90[6'h35:6'h35];
  assign T576 = T90[6'h36:6'h36];
  assign T577 = T90[6'h37:6'h37];
  assign T578 = T90[6'h38:6'h38];
  assign T579 = T90[6'h39:6'h39];
  assign T580 = T90[6'h3a:6'h3a];
  assign T581 = T90[6'h3b:6'h3b];
  assign T582 = T90[6'h3c:6'h3c];
  assign T583 = T90[6'h3d:6'h3d];
  assign T584 = T90[6'h3e:6'h3e];
  assign T585 = T90[6'h3f:6'h3f];
  assign T91 = T85 << 4'hc;
  assign T92 = T93 == 11'h0;
  assign T93 = R21[6'h3e:6'h34];
  assign T94 = T101 | T586;
  assign T586 = {2'h0, T95};
  assign T95 = T96 << 4'h9;
  assign T96 = T99 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T85 == 52'h0;
  assign T99 = T100 == 2'h3;
  assign T100 = T101[4'hb:4'ha];
  assign T101 = T108 + T587;
  assign T587 = {1'h0, T102};
  assign T102 = T107 ? 11'h0 : T103;
  assign T103 = 11'h400 | T588;
  assign T588 = {9'h0, T104};
  assign T104 = T105 ? 2'h2 : 2'h1;
  assign T105 = T92 & T106;
  assign T106 = T98 ^ 1'h1;
  assign T107 = T92 & T98;
  assign T108 = T92 ? T109 : T589;
  assign T589 = {1'h0, T93};
  assign T109 = T98 ? 12'h0 : T110;
  assign T110 = {6'h3f, T111};
  assign T111 = ~ T88;
  assign T112 = R21[6'h3f:6'h3f];
  assign T113 = {32'hffffffff, T114};
  assign T114 = {T144, T115};
  assign T115 = {T126, T116};
  assign T116 = T124 ? T118 : T117;
  assign T117 = R21[5'h16:1'h0];
  assign T118 = T119[5'h1e:4'h8];
  assign T119 = T123 << T120;
  assign T120 = ~ T590;
  assign T590 = T650 ? 5'h1f : T591;
  assign T591 = T649 ? 5'h1e : T592;
  assign T592 = T648 ? 5'h1d : T593;
  assign T593 = T647 ? 5'h1c : T594;
  assign T594 = T646 ? 5'h1b : T595;
  assign T595 = T645 ? 5'h1a : T596;
  assign T596 = T644 ? 5'h19 : T597;
  assign T597 = T643 ? 5'h18 : T598;
  assign T598 = T642 ? 5'h17 : T599;
  assign T599 = T641 ? 5'h16 : T600;
  assign T600 = T640 ? 5'h15 : T601;
  assign T601 = T639 ? 5'h14 : T602;
  assign T602 = T638 ? 5'h13 : T603;
  assign T603 = T637 ? 5'h12 : T604;
  assign T604 = T636 ? 5'h11 : T605;
  assign T605 = T635 ? 5'h10 : T606;
  assign T606 = T634 ? 4'hf : T607;
  assign T607 = T633 ? 4'he : T608;
  assign T608 = T632 ? 4'hd : T609;
  assign T609 = T631 ? 4'hc : T610;
  assign T610 = T630 ? 4'hb : T611;
  assign T611 = T629 ? 4'ha : T612;
  assign T612 = T628 ? 4'h9 : T613;
  assign T613 = T627 ? 4'h8 : T614;
  assign T614 = T626 ? 3'h7 : T615;
  assign T615 = T625 ? 3'h6 : T616;
  assign T616 = T624 ? 3'h5 : T617;
  assign T617 = T623 ? 3'h4 : T618;
  assign T618 = T622 ? 2'h3 : T619;
  assign T619 = T621 ? 2'h2 : T620;
  assign T620 = T122[1'h1:1'h1];
  assign T122 = T123[5'h1f:1'h0];
  assign T621 = T122[2'h2:2'h2];
  assign T622 = T122[2'h3:2'h3];
  assign T623 = T122[3'h4:3'h4];
  assign T624 = T122[3'h5:3'h5];
  assign T625 = T122[3'h6:3'h6];
  assign T626 = T122[3'h7:3'h7];
  assign T627 = T122[4'h8:4'h8];
  assign T628 = T122[4'h9:4'h9];
  assign T629 = T122[4'ha:4'ha];
  assign T630 = T122[4'hb:4'hb];
  assign T631 = T122[4'hc:4'hc];
  assign T632 = T122[4'hd:4'hd];
  assign T633 = T122[4'he:4'he];
  assign T634 = T122[4'hf:4'hf];
  assign T635 = T122[5'h10:5'h10];
  assign T636 = T122[5'h11:5'h11];
  assign T637 = T122[5'h12:5'h12];
  assign T638 = T122[5'h13:5'h13];
  assign T639 = T122[5'h14:5'h14];
  assign T640 = T122[5'h15:5'h15];
  assign T641 = T122[5'h16:5'h16];
  assign T642 = T122[5'h17:5'h17];
  assign T643 = T122[5'h18:5'h18];
  assign T644 = T122[5'h19:5'h19];
  assign T645 = T122[5'h1a:5'h1a];
  assign T646 = T122[5'h1b:5'h1b];
  assign T647 = T122[5'h1c:5'h1c];
  assign T648 = T122[5'h1d:5'h1d];
  assign T649 = T122[5'h1e:5'h1e];
  assign T650 = T122[5'h1f:5'h1f];
  assign T123 = T117 << 4'h9;
  assign T124 = T125 == 8'h0;
  assign T125 = R21[5'h1e:5'h17];
  assign T126 = T133 | T651;
  assign T651 = {2'h0, T127};
  assign T127 = T128 << 3'h6;
  assign T128 = T131 & T129;
  assign T129 = T130 ^ 1'h1;
  assign T130 = T117 == 23'h0;
  assign T131 = T132 == 2'h3;
  assign T132 = T133[4'h8:3'h7];
  assign T133 = T140 + T652;
  assign T652 = {1'h0, T134};
  assign T134 = T139 ? 8'h0 : T135;
  assign T135 = 8'h80 | T653;
  assign T653 = {6'h0, T136};
  assign T136 = T137 ? 2'h2 : 2'h1;
  assign T137 = T124 & T138;
  assign T138 = T130 ^ 1'h1;
  assign T139 = T124 & T130;
  assign T140 = T124 ? T141 : T654;
  assign T654 = {1'h0, T125};
  assign T141 = T130 ? 9'h0 : T142;
  assign T142 = {4'hf, T143};
  assign T143 = ~ T120;
  assign T144 = R21[5'h1f:5'h1f];
  assign T145 = {32'hffffffff, T146};
  assign T146 = {T24, T147};
  assign T147 = {T169, T148};
  assign T148 = T149[5'h16:1'h0];
  assign T149 = T153 ? T152 : T150;
  assign T150 = {1'h0, T151};
  assign T151 = T13[6'h3f:6'h28];
  assign T152 = T150 + 25'h1;
  assign T153 = T168 ? T163 : T154;
  assign T154 = T162 ? T161 : T155;
  assign T155 = T158 ? T156 : 1'h0;
  assign T156 = T157 & T8;
  assign T157 = T24 ^ 1'h1;
  assign T158 = R159 == 3'h3;
  assign T160 = io_in_valid ? io_in_bits_rm : R159;
  assign T161 = T24 & T8;
  assign T162 = R159 == 3'h2;
  assign T163 = T166 | T164;
  assign T164 = T165 == 2'h3;
  assign T165 = T10[1'h1:1'h0];
  assign T166 = T167 == 2'h3;
  assign T167 = T10[2'h2:1'h1];
  assign T168 = R159 == 3'h0;
  assign T169 = {T176, T170};
  assign T170 = T171[3'h7:1'h0];
  assign T171 = T173 + T655;
  assign T655 = {7'h0, T172};
  assign T172 = T149[5'h18:5'h18];
  assign T173 = {1'h0, T174};
  assign T174 = {1'h0, T175};
  assign T175 = ~ T14;
  assign T176 = T13[6'h3f:6'h3f];
  assign T177 = {T60, T178};
  assign T178 = {T198, T179};
  assign T179 = T180[6'h33:1'h0];
  assign T180 = T184 ? T183 : T181;
  assign T181 = {1'h0, T182};
  assign T182 = T51[6'h3f:4'hb];
  assign T183 = T181 + 54'h1;
  assign T184 = T197 ? T192 : T185;
  assign T185 = T191 ? T190 : T186;
  assign T186 = T189 ? T187 : 1'h0;
  assign T187 = T188 & T46;
  assign T188 = T60 ^ 1'h1;
  assign T189 = R159 == 3'h3;
  assign T190 = T60 & T46;
  assign T191 = R159 == 3'h2;
  assign T192 = T195 | T193;
  assign T193 = T194 == 2'h3;
  assign T194 = T48[1'h1:1'h0];
  assign T195 = T196 == 2'h3;
  assign T196 = T48[2'h2:1'h1];
  assign T197 = R159 == 3'h0;
  assign T198 = {T205, T199};
  assign T199 = T200[4'ha:1'h0];
  assign T200 = T202 + T656;
  assign T656 = {10'h0, T201};
  assign T201 = T180[6'h35:6'h35];
  assign T202 = {1'h0, T203};
  assign T203 = {4'h0, T204};
  assign T204 = ~ T52;
  assign T205 = T51[6'h3f:6'h3f];
  assign io_out_valid = R206;
  assign T657 = reset ? 1'h0 : R74;

  always @(posedge clk) begin
    if(R74) begin
      R0 <= R2;
    end
    if(R73) begin
      R2 <= mux_exc;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R29 <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      R38 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R42 <= io_in_bits_cmd;
    end
    if(reset) begin
      R73 <= 1'h0;
    end else begin
      R73 <= io_in_valid;
    end
    if(reset) begin
      R74 <= 1'h0;
    end else begin
      R74 <= R73;
    end
    if(R74) begin
      R75 <= R77;
    end
    if(R73) begin
      R77 <= mux_data;
    end
    if(io_in_valid) begin
      R159 <= io_in_bits_rm;
    end
    if(reset) begin
      R206 <= 1'h0;
    end else begin
      R206 <= R74;
    end
  end
endmodule

module FPToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc,
    input  io_lt
);

  reg [4:0] R0;
  wire[4:0] T1;
  wire[4:0] mux_exc;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] minmax_exc;
  wire T5;
  wire issnan2;
  wire T6;
  wire T7;
  wire T8;
  reg [64:0] R9;
  wire[64:0] T10;
  wire T11;
  reg  R12;
  wire T13;
  wire isnan2;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire issnan1;
  wire T18;
  wire T19;
  wire T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire T23;
  wire isnan1;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire isSgnj;
  wire[4:0] T28;
  reg [4:0] R29;
  wire[4:0] T30;
  wire[4:0] T31;
  wire[2:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[2:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire[11:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[1:0] T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire[27:0] T56;
  wire[51:0] T57;
  wire T58;
  wire[23:0] T59;
  wire[48:0] T60;
  wire[4:0] T61;
  wire[11:0] T62;
  wire[11:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire[48:0] T67;
  wire[47:0] T68;
  wire[23:0] T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[24:0] T76;
  wire[24:0] T77;
  wire[24:0] T78;
  wire[24:0] T79;
  wire[55:0] T80;
  wire[4:0] T81;
  wire[24:0] T82;
  wire[22:0] T83;
  wire[24:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  reg [2:0] R92;
  wire[2:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[1:0] T98;
  wire T99;
  wire[1:0] T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire[4:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[22:0] T115;
  wire T116;
  wire[2:0] T117;
  wire T118;
  wire T119;
  reg  R120;
  wire T200;
  reg [64:0] R121;
  wire[64:0] T122;
  wire[64:0] mux_data;
  wire[64:0] T123;
  wire[64:0] T124;
  wire[64:0] T125;
  wire[64:0] fsgnj;
  wire[32:0] T126;
  wire[31:0] T127;
  wire sign_s;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire sign_d;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire isLHS;
  wire T150;
  wire T151;
  wire T152;
  wire isMax;
  wire[64:0] T153;
  wire[32:0] T154;
  wire[31:0] T155;
  wire[22:0] T156;
  wire[22:0] T157;
  wire[22:0] T158;
  wire[22:0] T159;
  wire[22:0] T160;
  wire[22:0] T201;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[22:0] T170;
  wire[22:0] T202;
  wire[8:0] T171;
  wire[8:0] T172;
  wire[8:0] T173;
  wire[8:0] T174;
  wire[8:0] T175;
  wire[8:0] T176;
  wire[8:0] T177;
  wire T178;
  wire[8:0] T203;
  wire[6:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire[64:0] T182;
  wire[63:0] T183;
  wire[51:0] T184;
  wire[51:0] T185;
  wire[51:0] T186;
  wire[51:0] T204;
  wire[11:0] T187;
  wire[11:0] T188;
  wire[11:0] T189;
  wire[11:0] T190;
  wire T191;
  wire[11:0] T192;
  wire[7:0] T196;
  wire T193;
  wire[11:0] T205;
  wire[10:0] T194;
  wire T195;
  wire[11:0] T206;
  wire T197;
  wire T198;
  reg  R199;
  wire T207;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R9 = {3{$random}};
    R12 = {1{$random}};
    R21 = {3{$random}};
    R29 = {1{$random}};
    R92 = {1{$random}};
    R120 = {1{$random}};
    R121 = {3{$random}};
    R199 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R120 ? mux_exc : R0;
  assign mux_exc = T2;
  assign T2 = T118 ? T111 : T3;
  assign T3 = T108 ? T31 : T4;
  assign T4 = isSgnj ? 5'h0 : minmax_exc;
  assign minmax_exc = {T5, 4'h0};
  assign T5 = issnan1 | issnan2;
  assign issnan2 = isnan2 & T6;
  assign T6 = ~ T7;
  assign T7 = R12 ? T11 : T8;
  assign T8 = R9[6'h33:6'h33];
  assign T10 = io_in_valid ? io_in_bits_in2 : R9;
  assign T11 = R9[5'h16:5'h16];
  assign T13 = io_in_valid ? io_in_bits_single : R12;
  assign isnan2 = R12 ? T16 : T14;
  assign T14 = T15 == 3'h7;
  assign T15 = R9[6'h3f:6'h3d];
  assign T16 = T17 == 3'h7;
  assign T17 = R9[5'h1f:5'h1d];
  assign issnan1 = isnan1 & T18;
  assign T18 = ~ T19;
  assign T19 = R12 ? T23 : T20;
  assign T20 = R21[6'h33:6'h33];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = R21[5'h16:5'h16];
  assign isnan1 = R12 ? T26 : T24;
  assign T24 = T25 == 3'h7;
  assign T25 = R21[6'h3f:6'h3d];
  assign T26 = T27 == 3'h7;
  assign T27 = R21[5'h1f:5'h1d];
  assign isSgnj = T28 == 5'h4;
  assign T28 = R29 & 5'h5;
  assign T30 = io_in_valid ? io_in_bits_cmd : R29;
  assign T31 = {T103, T32};
  assign T32 = {T73, T33};
  assign T33 = {T71, T34};
  assign T34 = T45 | T35;
  assign T35 = T43 & T36;
  assign T36 = T37 ^ 1'h1;
  assign T37 = T41 | T38;
  assign T38 = T39 == 2'h3;
  assign T39 = T40[2'h2:1'h1];
  assign T40 = R21[6'h3f:6'h3d];
  assign T41 = T42 ^ 1'h1;
  assign T42 = T40 != 3'h0;
  assign T43 = T44 < 12'h76a;
  assign T44 = R21[6'h3f:6'h34];
  assign T45 = T49 | T46;
  assign T46 = T48 & T47;
  assign T47 = T37 ^ 1'h1;
  assign T48 = 12'h87f < T44;
  assign T49 = T51 & T50;
  assign T50 = T37 ^ 1'h1;
  assign T51 = T52 != 2'h0;
  assign T52 = T53[1'h1:1'h0];
  assign T53 = {T70, T54};
  assign T54 = T58 | T55;
  assign T55 = T56 != 28'h0;
  assign T56 = T57[5'h1b:1'h0];
  assign T57 = R21[6'h33:1'h0];
  assign T58 = T59 != 24'h0;
  assign T59 = T60[5'h17:1'h0];
  assign T60 = T67 >> T61;
  assign T61 = T62[3'h4:1'h0];
  assign T62 = T64 ? T63 : 12'h0;
  assign T63 = 12'h782 - T44;
  assign T64 = T66 & T65;
  assign T65 = T44 <= 12'h781;
  assign T66 = 12'h76a <= T44;
  assign T67 = {1'h1, T68};
  assign T68 = {T69, 24'h0};
  assign T69 = T57[6'h33:5'h1c];
  assign T70 = T60[5'h19:5'h18];
  assign T71 = T35 | T72;
  assign T72 = T64 & T49;
  assign T73 = T46 | T74;
  assign T74 = T102 & T75;
  assign T75 = T76[5'h18:5'h18];
  assign T76 = T85 ? T84 : T77;
  assign T77 = T82 | T78;
  assign T78 = ~ T79;
  assign T79 = T80[5'h18:1'h0];
  assign T80 = 25'h1ffffff << T81;
  assign T81 = T61;
  assign T82 = {2'h1, T83};
  assign T83 = T57[6'h33:5'h1d];
  assign T84 = T77 + 25'h1;
  assign T85 = T101 ? T96 : T86;
  assign T86 = T95 ? T94 : T87;
  assign T87 = T91 ? T88 : 1'h0;
  assign T88 = T89 & T49;
  assign T89 = T90 ^ 1'h1;
  assign T90 = R21[7'h40:7'h40];
  assign T91 = R92 == 3'h3;
  assign T93 = io_in_valid ? io_in_bits_rm : R92;
  assign T94 = T90 & T49;
  assign T95 = R92 == 3'h2;
  assign T96 = T99 | T97;
  assign T97 = T98 == 2'h3;
  assign T98 = T53[2'h2:1'h1];
  assign T99 = T100 == 2'h3;
  assign T100 = T53[1'h1:1'h0];
  assign T101 = R92 == 3'h0;
  assign T102 = T44 == 12'h87f;
  assign T103 = {T104, 1'h0};
  assign T104 = T107 & T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = T57[6'h33:6'h33];
  assign T107 = T40 == 3'h7;
  assign T108 = T109 & R12;
  assign T109 = T110 == 5'h0;
  assign T110 = R29 & 5'h4;
  assign T111 = T112 << 3'h4;
  assign T112 = T116 & T113;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115[5'h16:5'h16];
  assign T115 = R21[5'h16:1'h0];
  assign T116 = T117 == 3'h7;
  assign T117 = R21[5'h1f:5'h1d];
  assign T118 = T109 & T119;
  assign T119 = R12 ^ 1'h1;
  assign T200 = reset ? 1'h0 : io_in_valid;
  assign io_out_bits_data = R121;
  assign T122 = R120 ? mux_data : R121;
  assign mux_data = T123;
  assign T123 = T118 ? T182 : T124;
  assign T124 = T108 ? T153 : T125;
  assign T125 = T149 ? fsgnj : R9;
  assign fsgnj = {T137, T126};
  assign T126 = {sign_s, T127};
  assign T127 = R21[5'h1f:1'h0];
  assign sign_s = T131 ^ T128;
  assign T128 = T130 & T129;
  assign T129 = R9[6'h20:6'h20];
  assign T130 = R12 & isSgnj;
  assign T131 = T134 ? T133 : T132;
  assign T132 = R92[1'h0:1'h0];
  assign T133 = R21[6'h20:6'h20];
  assign T134 = T136 | T135;
  assign T135 = T130 ^ 1'h1;
  assign T136 = R92[1'h1:1'h1];
  assign T137 = {sign_d, T138};
  assign T138 = R21[6'h3f:6'h21];
  assign sign_d = T143 ^ T139;
  assign T139 = T141 & T140;
  assign T140 = R9[7'h40:7'h40];
  assign T141 = T142 & isSgnj;
  assign T142 = R12 ^ 1'h1;
  assign T143 = T146 ? T145 : T144;
  assign T144 = R92[1'h0:1'h0];
  assign T145 = R21[7'h40:7'h40];
  assign T146 = T148 | T147;
  assign T147 = T141 ^ 1'h1;
  assign T148 = R92[1'h1:1'h1];
  assign T149 = isSgnj | isLHS;
  assign isLHS = isnan2 | T150;
  assign T150 = T152 & T151;
  assign T151 = isnan1 ^ 1'h1;
  assign T152 = isMax != io_lt;
  assign isMax = R92[1'h0:1'h0];
  assign T153 = {32'hffffffff, T154};
  assign T154 = {T90, T155};
  assign T155 = {T171, T156};
  assign T156 = T37 ? T170 : T157;
  assign T157 = T46 ? T160 : T158;
  assign T158 = T35 ? 23'h0 : T159;
  assign T159 = T76[5'h16:1'h0];
  assign T160 = 23'h0 - T201;
  assign T201 = {22'h0, T161};
  assign T161 = T162 ^ 1'h1;
  assign T162 = T164 | T163;
  assign T163 = R92 == 3'h0;
  assign T164 = T168 | T165;
  assign T165 = T167 & T166;
  assign T166 = T90 ^ 1'h1;
  assign T167 = R92 == 3'h3;
  assign T168 = T169 & T90;
  assign T169 = R92 == 3'h2;
  assign T170 = 23'h0 - T202;
  assign T202 = {22'h0, T107};
  assign T171 = T37 ? T181 : T172;
  assign T172 = T46 ? T180 : T173;
  assign T173 = T35 ? T203 : T174;
  assign T174 = T178 ? T177 : T175;
  assign T175 = T176 + 9'h100;
  assign T176 = T44[4'h8:1'h0];
  assign T177 = T175 + 9'h1;
  assign T178 = T76[5'h18:5'h18];
  assign T203 = {2'h0, T179};
  assign T179 = T164 ? 7'h6b : 7'h0;
  assign T180 = T162 ? 9'h180 : 9'h17f;
  assign T181 = T40 << 3'h6;
  assign T182 = {T198, T183};
  assign T183 = {T187, T184};
  assign T184 = T186 | T185;
  assign T185 = T115 << 5'h1d;
  assign T186 = 52'h0 - T204;
  assign T204 = {51'h0, T116};
  assign T187 = T197 ? T206 : T188;
  assign T188 = T195 ? T205 : T189;
  assign T189 = T193 ? T192 : T190;
  assign T190 = T191 ? 12'hc00 : 12'he00;
  assign T191 = T117 < 3'h7;
  assign T192 = {4'h8, T196};
  assign T196 = R21[5'h1e:5'h17];
  assign T193 = T117 < 3'h6;
  assign T205 = {1'h0, T194};
  assign T194 = {3'h7, T196};
  assign T195 = T117 < 3'h4;
  assign T206 = {4'h0, T196};
  assign T197 = T117 < 3'h1;
  assign T198 = R21[6'h20:6'h20];
  assign io_out_valid = R199;
  assign T207 = reset ? 1'h0 : R120;

  always @(posedge clk) begin
    if(R120) begin
      R0 <= mux_exc;
    end
    if(io_in_valid) begin
      R9 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      R12 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R29 <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      R92 <= io_in_bits_rm;
    end
    if(reset) begin
      R120 <= 1'h0;
    end else begin
      R120 <= io_in_valid;
    end
    if(R120) begin
      R121 <= mux_data;
    end
    if(reset) begin
      R199 <= 1'h0;
    end else begin
      R199 <= R120;
    end
  end
endmodule

module FPU(input clk, input reset,
    input  io_ctrl_valid,
    output io_ctrl_fcsr_rdy,
    output io_ctrl_nack_mem,
    output io_ctrl_illegal_rm,
    input  io_ctrl_killx,
    input  io_ctrl_killm,
    output[4:0] io_ctrl_dec_cmd,
    output io_ctrl_dec_ldst,
    output io_ctrl_dec_wen,
    output io_ctrl_dec_ren1,
    output io_ctrl_dec_ren2,
    output io_ctrl_dec_ren3,
    output io_ctrl_dec_swap23,
    output io_ctrl_dec_single,
    output io_ctrl_dec_fromint,
    output io_ctrl_dec_toint,
    output io_ctrl_dec_fastpipe,
    output io_ctrl_dec_fma,
    output io_ctrl_dec_round,
    output io_ctrl_sboard_set,
    output io_ctrl_sboard_clr,
    output[4:0] io_ctrl_sboard_clra,
    input [31:0] io_dpath_inst,
    input [63:0] io_dpath_fromint_data,
    input [2:0] io_dpath_fcsr_rm,
    output io_dpath_fcsr_flags_valid,
    output[4:0] io_dpath_fcsr_flags_bits,
    output[63:0] io_dpath_store_data,
    output[63:0] io_dpath_toint_data,
    input  io_dpath_dmem_resp_val,
    input [2:0] io_dpath_dmem_resp_type,
    input [4:0] io_dpath_dmem_resp_tag,
    input [63:0] io_dpath_dmem_resp_data
);

  wire[64:0] req_in3;
  wire[64:0] ex_rs3;
  reg [64:0] regfile [31:0];
  wire[64:0] T0;
  wire[64:0] T223;
  wire[96:0] wdata;
  wire[96:0] T224;
  wire[64:0] T1;
  wire T2;
  wire[1:0] T3;
  wire[1:0] wsrc;
  reg [6:0] winfo_0;
  wire[6:0] T4;
  wire[6:0] T5;
  reg [6:0] winfo_1;
  wire[6:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] memLatencyMask;
  wire[1:0] T10;
  wire T11;
  wire T12;
  reg  mem_ctrl_single;
  wire T13;
  reg  ex_ctrl_single;
  wire T14;
  reg  ex_reg_valid;
  wire T225;
  reg  mem_ctrl_fma;
  wire T15;
  reg  ex_ctrl_fma;
  wire T16;
  wire[1:0] T17;
  wire[1:0] T226;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  reg  mem_ctrl_fromint;
  wire T21;
  reg  ex_ctrl_fromint;
  wire T22;
  wire[1:0] T227;
  reg  mem_ctrl_fastpipe;
  wire T23;
  reg  ex_ctrl_fastpipe;
  wire T24;
  wire T25;
  reg  write_port_busy;
  wire T26;
  wire T27;
  wire T28;
  wire[3:0] T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire T32;
  wire T33;
  wire[3:0] T34;
  wire[3:0] T228;
  wire[2:0] T35;
  wire T36;
  wire[3:0] T37;
  wire[3:0] T38;
  wire[3:0] T229;
  wire[2:0] T39;
  wire[3:0] T230;
  reg [1:0] wen;
  wire[1:0] T231;
  wire[1:0] T40;
  wire[1:0] T232;
  wire T41;
  wire[1:0] T42;
  wire[1:0] T233;
  wire T43;
  wire T44;
  wire T45;
  wire killm;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire[2:0] T50;
  wire T51;
  wire T52;
  wire[2:0] T53;
  wire[2:0] T234;
  wire[1:0] T54;
  wire T55;
  wire[2:0] T56;
  wire[2:0] T57;
  wire[2:0] T235;
  wire[1:0] T58;
  wire[2:0] T236;
  wire mem_wen;
  wire T59;
  wire T60;
  reg  mem_reg_valid;
  wire T237;
  wire T61;
  wire T62;
  wire T63;
  wire[6:0] mem_winfo;
  wire[4:0] T64;
  reg [31:0] mem_reg_inst;
  wire[31:0] T65;
  reg [31:0] ex_reg_inst;
  wire[31:0] T66;
  wire[1:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire T73;
  wire[1:0] T238;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire[96:0] T79;
  wire[96:0] T80;
  wire[96:0] T239;
  wire T81;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire[4:0] waddr;
  wire[4:0] T85;
  wire[64:0] T86;
  wire[64:0] load_wb_data_recoded;
  wire[64:0] rec_d;
  wire[63:0] T87;
  wire[51:0] T88;
  wire[51:0] T89;
  reg [63:0] load_wb_data;
  wire[63:0] T90;
  wire[51:0] T91;
  wire[126:0] T92;
  wire[5:0] T93;
  wire[5:0] T240;
  wire[5:0] T241;
  wire[5:0] T242;
  wire[5:0] T243;
  wire[5:0] T244;
  wire[5:0] T245;
  wire[5:0] T246;
  wire[5:0] T247;
  wire[5:0] T248;
  wire[5:0] T249;
  wire[5:0] T250;
  wire[5:0] T251;
  wire[5:0] T252;
  wire[5:0] T253;
  wire[5:0] T254;
  wire[5:0] T255;
  wire[5:0] T256;
  wire[5:0] T257;
  wire[5:0] T258;
  wire[5:0] T259;
  wire[5:0] T260;
  wire[5:0] T261;
  wire[5:0] T262;
  wire[5:0] T263;
  wire[5:0] T264;
  wire[5:0] T265;
  wire[5:0] T266;
  wire[5:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[5:0] T270;
  wire[5:0] T271;
  wire[4:0] T272;
  wire[4:0] T273;
  wire[4:0] T274;
  wire[4:0] T275;
  wire[4:0] T276;
  wire[4:0] T277;
  wire[4:0] T278;
  wire[4:0] T279;
  wire[4:0] T280;
  wire[4:0] T281;
  wire[4:0] T282;
  wire[4:0] T283;
  wire[4:0] T284;
  wire[4:0] T285;
  wire[4:0] T286;
  wire[4:0] T287;
  wire[3:0] T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[3:0] T294;
  wire[3:0] T295;
  wire[2:0] T296;
  wire[2:0] T297;
  wire[2:0] T298;
  wire[2:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire T302;
  wire[63:0] T95;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire[63:0] T96;
  wire T97;
  wire[10:0] T98;
  wire[11:0] T99;
  wire[11:0] T365;
  wire[9:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire[1:0] T105;
  wire[11:0] T106;
  wire[11:0] T366;
  wire[10:0] T107;
  wire[10:0] T108;
  wire[10:0] T367;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[11:0] T113;
  wire[11:0] T368;
  wire[11:0] T114;
  wire[11:0] T115;
  wire[5:0] T116;
  wire T117;
  wire[64:0] T118;
  wire[32:0] rec_s;
  wire[31:0] T119;
  wire[22:0] T120;
  wire[22:0] T121;
  wire[22:0] T122;
  wire[62:0] T123;
  wire[4:0] T124;
  wire[4:0] T369;
  wire[4:0] T370;
  wire[4:0] T371;
  wire[4:0] T372;
  wire[4:0] T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire[4:0] T377;
  wire[4:0] T378;
  wire[4:0] T379;
  wire[4:0] T380;
  wire[4:0] T381;
  wire[4:0] T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[3:0] T390;
  wire[3:0] T391;
  wire[3:0] T392;
  wire[2:0] T393;
  wire[2:0] T394;
  wire[2:0] T395;
  wire[2:0] T396;
  wire[1:0] T397;
  wire[1:0] T398;
  wire T399;
  wire[31:0] T126;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire[31:0] T127;
  wire T128;
  wire[7:0] T129;
  wire[8:0] T130;
  wire[8:0] T430;
  wire[6:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[1:0] T136;
  wire[8:0] T137;
  wire[8:0] T431;
  wire[7:0] T138;
  wire[7:0] T139;
  wire[7:0] T432;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[8:0] T144;
  wire[8:0] T433;
  wire[8:0] T145;
  wire[8:0] T146;
  wire[4:0] T147;
  wire T148;
  reg  load_wb_single;
  wire T149;
  wire T150;
  wire T151;
  wire[3:0] T434;
  wire T152;
  wire[3:0] T435;
  reg  load_wb;
  reg [4:0] load_wb_tag;
  wire[4:0] T153;
  reg [4:0] ex_ra3;
  wire[4:0] T154;
  wire[4:0] T155;
  wire[4:0] T156;
  wire T157;
  wire[4:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[64:0] req_in2;
  wire[64:0] ex_rs2;
  reg [4:0] ex_ra2;
  wire[4:0] T163;
  wire[4:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[64:0] req_in1;
  wire[64:0] ex_rs1;
  reg [4:0] ex_ra1;
  wire[4:0] T169;
  wire[4:0] T170;
  wire[4:0] T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire[1:0] req_typ;
  wire[1:0] T175;
  wire[2:0] req_rm;
  wire[2:0] ex_rm;
  wire[2:0] T176;
  wire T177;
  wire[2:0] T178;
  wire req_round;
  reg  ex_ctrl_round;
  wire T179;
  wire req_fma;
  wire req_fastpipe;
  wire req_toint;
  reg  ex_ctrl_toint;
  wire T180;
  wire req_fromint;
  wire req_single;
  wire req_swap23;
  reg  ex_ctrl_swap23;
  wire T181;
  wire req_ren3;
  reg  ex_ctrl_ren3;
  wire T182;
  wire req_ren2;
  reg  ex_ctrl_ren2;
  wire T183;
  wire req_ren1;
  reg  ex_ctrl_ren1;
  wire T184;
  wire req_wen;
  reg  ex_ctrl_wen;
  wire T185;
  wire req_ldst;
  reg  ex_ctrl_ldst;
  wire T186;
  wire[4:0] req_cmd;
  reg [4:0] ex_ctrl_cmd;
  wire[4:0] T187;
  wire T188;
  wire[64:0] T436;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire[4:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire[4:0] T199;
  wire[4:0] T200;
  wire[4:0] wexc;
  wire[4:0] T201;
  wire T202;
  wire[1:0] T203;
  wire[4:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire[4:0] T208;
  reg [4:0] wb_toint_exc;
  wire[4:0] T209;
  reg  mem_ctrl_toint;
  wire T210;
  wire wb_toint_valid;
  reg  wb_ctrl_toint;
  wire T211;
  reg  wb_reg_valid;
  wire T437;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  reg  R217;
  wire T218;
  wire T219;
  wire T220;
  wire fp_inflight;
  wire T221;
  wire T222;
  wire[4:0] fp_decoder_io_sigs_cmd;
  wire fp_decoder_io_sigs_ldst;
  wire fp_decoder_io_sigs_wen;
  wire fp_decoder_io_sigs_ren1;
  wire fp_decoder_io_sigs_ren2;
  wire fp_decoder_io_sigs_ren3;
  wire fp_decoder_io_sigs_swap23;
  wire fp_decoder_io_sigs_single;
  wire fp_decoder_io_sigs_fromint;
  wire fp_decoder_io_sigs_toint;
  wire fp_decoder_io_sigs_fastpipe;
  wire fp_decoder_io_sigs_fma;
  wire fp_decoder_io_sigs_round;
  wire[64:0] ifpu_io_out_bits_data;
  wire[4:0] ifpu_io_out_bits_exc;
  wire[64:0] fpmu_io_out_bits_data;
  wire[4:0] fpmu_io_out_bits_exc;
  wire[64:0] sfma_io_out_bits_data;
  wire[4:0] sfma_io_out_bits_exc;
  wire[64:0] dfma_io_out_bits_data;
  wire[4:0] dfma_io_out_bits_exc;
  wire fpiu_io_out_bits_lt;
  wire[63:0] fpiu_io_out_bits_store;
  wire[63:0] fpiu_io_out_bits_toint;
  wire[4:0] fpiu_io_out_bits_exc;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 32; initvar = initvar+1)
      regfile[initvar] = {3{$random}};
    winfo_0 = {1{$random}};
    winfo_1 = {1{$random}};
    mem_ctrl_single = {1{$random}};
    ex_ctrl_single = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_ctrl_fma = {1{$random}};
    ex_ctrl_fma = {1{$random}};
    mem_ctrl_fromint = {1{$random}};
    ex_ctrl_fromint = {1{$random}};
    mem_ctrl_fastpipe = {1{$random}};
    ex_ctrl_fastpipe = {1{$random}};
    write_port_busy = {1{$random}};
    wen = {1{$random}};
    mem_reg_valid = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    load_wb_data = {2{$random}};
    load_wb_single = {1{$random}};
    load_wb = {1{$random}};
    load_wb_tag = {1{$random}};
    ex_ra3 = {1{$random}};
    ex_ra2 = {1{$random}};
    ex_ra1 = {1{$random}};
    ex_ctrl_round = {1{$random}};
    ex_ctrl_toint = {1{$random}};
    ex_ctrl_swap23 = {1{$random}};
    ex_ctrl_ren3 = {1{$random}};
    ex_ctrl_ren2 = {1{$random}};
    ex_ctrl_ren1 = {1{$random}};
    ex_ctrl_wen = {1{$random}};
    ex_ctrl_ldst = {1{$random}};
    ex_ctrl_cmd = {1{$random}};
    wb_toint_exc = {1{$random}};
    mem_ctrl_toint = {1{$random}};
    wb_ctrl_toint = {1{$random}};
    wb_reg_valid = {1{$random}};
    R217 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign req_in3 = ex_rs3;
  assign ex_rs3 = regfile[ex_ra3];
  assign T223 = wdata[7'h40:1'h0];
  assign wdata = T82 ? T79 : T224;
  assign T224 = {32'h0, T1};
  assign T1 = T2 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data;
  assign T2 = T3[1'h0:1'h0];
  assign T3 = wsrc;
  assign wsrc = winfo_0 >> 3'h5;
  assign T4 = T75 ? mem_winfo : T5;
  assign T5 = T63 ? winfo_1 : winfo_0;
  assign T6 = T7 ? mem_winfo : winfo_1;
  assign T7 = mem_wen & T8;
  assign T8 = T25 & T9;
  assign T9 = memLatencyMask[1'h1:1'h1];
  assign memLatencyMask = T17 | T10;
  assign T10 = T11 ? 2'h2 : 2'h0;
  assign T11 = mem_ctrl_fma & T12;
  assign T12 = mem_ctrl_single ^ 1'h1;
  assign T13 = ex_reg_valid ? ex_ctrl_single : mem_ctrl_single;
  assign T14 = io_ctrl_valid ? fp_decoder_io_sigs_single : ex_ctrl_single;
  assign T225 = reset ? 1'h0 : io_ctrl_valid;
  assign T15 = ex_reg_valid ? ex_ctrl_fma : mem_ctrl_fma;
  assign T16 = io_ctrl_valid ? fp_decoder_io_sigs_fma : ex_ctrl_fma;
  assign T17 = T19 | T226;
  assign T226 = {1'h0, T18};
  assign T18 = mem_ctrl_fma & mem_ctrl_single;
  assign T19 = T227 | T20;
  assign T20 = mem_ctrl_fromint ? 2'h2 : 2'h0;
  assign T21 = ex_reg_valid ? ex_ctrl_fromint : mem_ctrl_fromint;
  assign T22 = io_ctrl_valid ? fp_decoder_io_sigs_fromint : ex_ctrl_fromint;
  assign T227 = {1'h0, mem_ctrl_fastpipe};
  assign T23 = ex_reg_valid ? ex_ctrl_fastpipe : mem_ctrl_fastpipe;
  assign T24 = io_ctrl_valid ? fp_decoder_io_sigs_fastpipe : ex_ctrl_fastpipe;
  assign T25 = write_port_busy ^ 1'h1;
  assign T26 = ex_reg_valid ? T27 : write_port_busy;
  assign T27 = T46 | T28;
  assign T28 = T29 != 4'h0;
  assign T29 = T230 & T30;
  assign T30 = T34 | T31;
  assign T31 = T32 ? 4'h8 : 4'h0;
  assign T32 = ex_ctrl_fma & T33;
  assign T33 = ex_ctrl_single ^ 1'h1;
  assign T34 = T37 | T228;
  assign T228 = {1'h0, T35};
  assign T35 = T36 ? 3'h4 : 3'h0;
  assign T36 = ex_ctrl_fma & ex_ctrl_single;
  assign T37 = T229 | T38;
  assign T38 = ex_ctrl_fromint ? 4'h8 : 4'h0;
  assign T229 = {1'h0, T39};
  assign T39 = ex_ctrl_fastpipe ? 3'h4 : 3'h0;
  assign T230 = {2'h0, wen};
  assign T231 = reset ? 2'h0 : T40;
  assign T40 = T44 ? T42 : T232;
  assign T232 = {1'h0, T41};
  assign T41 = wen >> 1'h1;
  assign T42 = T233 | memLatencyMask;
  assign T233 = {1'h0, T43};
  assign T43 = wen >> 1'h1;
  assign T44 = mem_wen & T45;
  assign T45 = killm ^ 1'h1;
  assign killm = io_ctrl_killm | io_ctrl_nack_mem;
  assign T46 = mem_wen & T47;
  assign T47 = T48 != 3'h0;
  assign T48 = T236 & T49;
  assign T49 = T53 | T50;
  assign T50 = T51 ? 3'h4 : 3'h0;
  assign T51 = ex_ctrl_fma & T52;
  assign T52 = ex_ctrl_single ^ 1'h1;
  assign T53 = T56 | T234;
  assign T234 = {1'h0, T54};
  assign T54 = T55 ? 2'h2 : 2'h0;
  assign T55 = ex_ctrl_fma & ex_ctrl_single;
  assign T56 = T235 | T57;
  assign T57 = ex_ctrl_fromint ? 3'h4 : 3'h0;
  assign T235 = {1'h0, T58};
  assign T58 = ex_ctrl_fastpipe ? 2'h2 : 2'h0;
  assign T236 = {1'h0, memLatencyMask};
  assign mem_wen = mem_reg_valid & T59;
  assign T59 = T60 | mem_ctrl_fromint;
  assign T60 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T237 = reset ? 1'h0 : T61;
  assign T61 = ex_reg_valid & T62;
  assign T62 = io_ctrl_killx ^ 1'h1;
  assign T63 = wen[1'h1:1'h1];
  assign mem_winfo = {T67, T64};
  assign T64 = mem_reg_inst[4'hb:3'h7];
  assign T65 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T66 = io_ctrl_valid ? io_dpath_inst : ex_reg_inst;
  assign T67 = T71 | T68;
  assign T68 = T69 ? 2'h3 : 2'h0;
  assign T69 = mem_ctrl_fma & T70;
  assign T70 = mem_ctrl_single ^ 1'h1;
  assign T71 = T238 | T72;
  assign T72 = T73 ? 2'h2 : 2'h0;
  assign T73 = mem_ctrl_fma & mem_ctrl_single;
  assign T238 = {1'h0, T74};
  assign T74 = 1'h0 | mem_ctrl_fromint;
  assign T75 = mem_wen & T76;
  assign T76 = T78 & T77;
  assign T77 = memLatencyMask[1'h0:1'h0];
  assign T78 = write_port_busy ^ 1'h1;
  assign T79 = T81 ? T239 : T80;
  assign T80 = {32'hffffffff, sfma_io_out_bits_data};
  assign T239 = {32'h0, dfma_io_out_bits_data};
  assign T81 = T3[1'h0:1'h0];
  assign T82 = T3[1'h1:1'h1];
  assign T83 = wen[1'h0:1'h0];
  assign T84 = waddr[3'h4:1'h0];
  assign waddr = T85;
  assign T85 = winfo_0[3'h4:1'h0];
  assign load_wb_data_recoded = load_wb_single ? T118 : rec_d;
  assign rec_d = {T117, T87};
  assign T87 = {T99, T88};
  assign T88 = T97 ? T91 : T89;
  assign T89 = load_wb_data[6'h33:1'h0];
  assign T90 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_data : load_wb_data;
  assign T91 = T92[6'h3e:4'hb];
  assign T92 = T96 << T93;
  assign T93 = ~ T240;
  assign T240 = T364 ? 6'h3f : T241;
  assign T241 = T363 ? 6'h3e : T242;
  assign T242 = T362 ? 6'h3d : T243;
  assign T243 = T361 ? 6'h3c : T244;
  assign T244 = T360 ? 6'h3b : T245;
  assign T245 = T359 ? 6'h3a : T246;
  assign T246 = T358 ? 6'h39 : T247;
  assign T247 = T357 ? 6'h38 : T248;
  assign T248 = T356 ? 6'h37 : T249;
  assign T249 = T355 ? 6'h36 : T250;
  assign T250 = T354 ? 6'h35 : T251;
  assign T251 = T353 ? 6'h34 : T252;
  assign T252 = T352 ? 6'h33 : T253;
  assign T253 = T351 ? 6'h32 : T254;
  assign T254 = T350 ? 6'h31 : T255;
  assign T255 = T349 ? 6'h30 : T256;
  assign T256 = T348 ? 6'h2f : T257;
  assign T257 = T347 ? 6'h2e : T258;
  assign T258 = T346 ? 6'h2d : T259;
  assign T259 = T345 ? 6'h2c : T260;
  assign T260 = T344 ? 6'h2b : T261;
  assign T261 = T343 ? 6'h2a : T262;
  assign T262 = T342 ? 6'h29 : T263;
  assign T263 = T341 ? 6'h28 : T264;
  assign T264 = T340 ? 6'h27 : T265;
  assign T265 = T339 ? 6'h26 : T266;
  assign T266 = T338 ? 6'h25 : T267;
  assign T267 = T337 ? 6'h24 : T268;
  assign T268 = T336 ? 6'h23 : T269;
  assign T269 = T335 ? 6'h22 : T270;
  assign T270 = T334 ? 6'h21 : T271;
  assign T271 = T333 ? 6'h20 : T272;
  assign T272 = T332 ? 5'h1f : T273;
  assign T273 = T331 ? 5'h1e : T274;
  assign T274 = T330 ? 5'h1d : T275;
  assign T275 = T329 ? 5'h1c : T276;
  assign T276 = T328 ? 5'h1b : T277;
  assign T277 = T327 ? 5'h1a : T278;
  assign T278 = T326 ? 5'h19 : T279;
  assign T279 = T325 ? 5'h18 : T280;
  assign T280 = T324 ? 5'h17 : T281;
  assign T281 = T323 ? 5'h16 : T282;
  assign T282 = T322 ? 5'h15 : T283;
  assign T283 = T321 ? 5'h14 : T284;
  assign T284 = T320 ? 5'h13 : T285;
  assign T285 = T319 ? 5'h12 : T286;
  assign T286 = T318 ? 5'h11 : T287;
  assign T287 = T317 ? 5'h10 : T288;
  assign T288 = T316 ? 4'hf : T289;
  assign T289 = T315 ? 4'he : T290;
  assign T290 = T314 ? 4'hd : T291;
  assign T291 = T313 ? 4'hc : T292;
  assign T292 = T312 ? 4'hb : T293;
  assign T293 = T311 ? 4'ha : T294;
  assign T294 = T310 ? 4'h9 : T295;
  assign T295 = T309 ? 4'h8 : T296;
  assign T296 = T308 ? 3'h7 : T297;
  assign T297 = T307 ? 3'h6 : T298;
  assign T298 = T306 ? 3'h5 : T299;
  assign T299 = T305 ? 3'h4 : T300;
  assign T300 = T304 ? 2'h3 : T301;
  assign T301 = T303 ? 2'h2 : T302;
  assign T302 = T95[1'h1:1'h1];
  assign T95 = T96[6'h3f:1'h0];
  assign T303 = T95[2'h2:2'h2];
  assign T304 = T95[2'h3:2'h3];
  assign T305 = T95[3'h4:3'h4];
  assign T306 = T95[3'h5:3'h5];
  assign T307 = T95[3'h6:3'h6];
  assign T308 = T95[3'h7:3'h7];
  assign T309 = T95[4'h8:4'h8];
  assign T310 = T95[4'h9:4'h9];
  assign T311 = T95[4'ha:4'ha];
  assign T312 = T95[4'hb:4'hb];
  assign T313 = T95[4'hc:4'hc];
  assign T314 = T95[4'hd:4'hd];
  assign T315 = T95[4'he:4'he];
  assign T316 = T95[4'hf:4'hf];
  assign T317 = T95[5'h10:5'h10];
  assign T318 = T95[5'h11:5'h11];
  assign T319 = T95[5'h12:5'h12];
  assign T320 = T95[5'h13:5'h13];
  assign T321 = T95[5'h14:5'h14];
  assign T322 = T95[5'h15:5'h15];
  assign T323 = T95[5'h16:5'h16];
  assign T324 = T95[5'h17:5'h17];
  assign T325 = T95[5'h18:5'h18];
  assign T326 = T95[5'h19:5'h19];
  assign T327 = T95[5'h1a:5'h1a];
  assign T328 = T95[5'h1b:5'h1b];
  assign T329 = T95[5'h1c:5'h1c];
  assign T330 = T95[5'h1d:5'h1d];
  assign T331 = T95[5'h1e:5'h1e];
  assign T332 = T95[5'h1f:5'h1f];
  assign T333 = T95[6'h20:6'h20];
  assign T334 = T95[6'h21:6'h21];
  assign T335 = T95[6'h22:6'h22];
  assign T336 = T95[6'h23:6'h23];
  assign T337 = T95[6'h24:6'h24];
  assign T338 = T95[6'h25:6'h25];
  assign T339 = T95[6'h26:6'h26];
  assign T340 = T95[6'h27:6'h27];
  assign T341 = T95[6'h28:6'h28];
  assign T342 = T95[6'h29:6'h29];
  assign T343 = T95[6'h2a:6'h2a];
  assign T344 = T95[6'h2b:6'h2b];
  assign T345 = T95[6'h2c:6'h2c];
  assign T346 = T95[6'h2d:6'h2d];
  assign T347 = T95[6'h2e:6'h2e];
  assign T348 = T95[6'h2f:6'h2f];
  assign T349 = T95[6'h30:6'h30];
  assign T350 = T95[6'h31:6'h31];
  assign T351 = T95[6'h32:6'h32];
  assign T352 = T95[6'h33:6'h33];
  assign T353 = T95[6'h34:6'h34];
  assign T354 = T95[6'h35:6'h35];
  assign T355 = T95[6'h36:6'h36];
  assign T356 = T95[6'h37:6'h37];
  assign T357 = T95[6'h38:6'h38];
  assign T358 = T95[6'h39:6'h39];
  assign T359 = T95[6'h3a:6'h3a];
  assign T360 = T95[6'h3b:6'h3b];
  assign T361 = T95[6'h3c:6'h3c];
  assign T362 = T95[6'h3d:6'h3d];
  assign T363 = T95[6'h3e:6'h3e];
  assign T364 = T95[6'h3f:6'h3f];
  assign T96 = T89 << 4'hc;
  assign T97 = T98 == 11'h0;
  assign T98 = load_wb_data[6'h3e:6'h34];
  assign T99 = T106 | T365;
  assign T365 = {2'h0, T100};
  assign T100 = T101 << 4'h9;
  assign T101 = T104 & T102;
  assign T102 = T103 ^ 1'h1;
  assign T103 = T89 == 52'h0;
  assign T104 = T105 == 2'h3;
  assign T105 = T106[4'hb:4'ha];
  assign T106 = T113 + T366;
  assign T366 = {1'h0, T107};
  assign T107 = T112 ? 11'h0 : T108;
  assign T108 = 11'h400 | T367;
  assign T367 = {9'h0, T109};
  assign T109 = T110 ? 2'h2 : 2'h1;
  assign T110 = T97 & T111;
  assign T111 = T103 ^ 1'h1;
  assign T112 = T97 & T103;
  assign T113 = T97 ? T114 : T368;
  assign T368 = {1'h0, T98};
  assign T114 = T103 ? 12'h0 : T115;
  assign T115 = {6'h3f, T116};
  assign T116 = ~ T93;
  assign T117 = load_wb_data[6'h3f:6'h3f];
  assign T118 = {32'hffffffff, rec_s};
  assign rec_s = {T148, T119};
  assign T119 = {T130, T120};
  assign T120 = T128 ? T122 : T121;
  assign T121 = load_wb_data[5'h16:1'h0];
  assign T122 = T123[5'h1e:4'h8];
  assign T123 = T127 << T124;
  assign T124 = ~ T369;
  assign T369 = T429 ? 5'h1f : T370;
  assign T370 = T428 ? 5'h1e : T371;
  assign T371 = T427 ? 5'h1d : T372;
  assign T372 = T426 ? 5'h1c : T373;
  assign T373 = T425 ? 5'h1b : T374;
  assign T374 = T424 ? 5'h1a : T375;
  assign T375 = T423 ? 5'h19 : T376;
  assign T376 = T422 ? 5'h18 : T377;
  assign T377 = T421 ? 5'h17 : T378;
  assign T378 = T420 ? 5'h16 : T379;
  assign T379 = T419 ? 5'h15 : T380;
  assign T380 = T418 ? 5'h14 : T381;
  assign T381 = T417 ? 5'h13 : T382;
  assign T382 = T416 ? 5'h12 : T383;
  assign T383 = T415 ? 5'h11 : T384;
  assign T384 = T414 ? 5'h10 : T385;
  assign T385 = T413 ? 4'hf : T386;
  assign T386 = T412 ? 4'he : T387;
  assign T387 = T411 ? 4'hd : T388;
  assign T388 = T410 ? 4'hc : T389;
  assign T389 = T409 ? 4'hb : T390;
  assign T390 = T408 ? 4'ha : T391;
  assign T391 = T407 ? 4'h9 : T392;
  assign T392 = T406 ? 4'h8 : T393;
  assign T393 = T405 ? 3'h7 : T394;
  assign T394 = T404 ? 3'h6 : T395;
  assign T395 = T403 ? 3'h5 : T396;
  assign T396 = T402 ? 3'h4 : T397;
  assign T397 = T401 ? 2'h3 : T398;
  assign T398 = T400 ? 2'h2 : T399;
  assign T399 = T126[1'h1:1'h1];
  assign T126 = T127[5'h1f:1'h0];
  assign T400 = T126[2'h2:2'h2];
  assign T401 = T126[2'h3:2'h3];
  assign T402 = T126[3'h4:3'h4];
  assign T403 = T126[3'h5:3'h5];
  assign T404 = T126[3'h6:3'h6];
  assign T405 = T126[3'h7:3'h7];
  assign T406 = T126[4'h8:4'h8];
  assign T407 = T126[4'h9:4'h9];
  assign T408 = T126[4'ha:4'ha];
  assign T409 = T126[4'hb:4'hb];
  assign T410 = T126[4'hc:4'hc];
  assign T411 = T126[4'hd:4'hd];
  assign T412 = T126[4'he:4'he];
  assign T413 = T126[4'hf:4'hf];
  assign T414 = T126[5'h10:5'h10];
  assign T415 = T126[5'h11:5'h11];
  assign T416 = T126[5'h12:5'h12];
  assign T417 = T126[5'h13:5'h13];
  assign T418 = T126[5'h14:5'h14];
  assign T419 = T126[5'h15:5'h15];
  assign T420 = T126[5'h16:5'h16];
  assign T421 = T126[5'h17:5'h17];
  assign T422 = T126[5'h18:5'h18];
  assign T423 = T126[5'h19:5'h19];
  assign T424 = T126[5'h1a:5'h1a];
  assign T425 = T126[5'h1b:5'h1b];
  assign T426 = T126[5'h1c:5'h1c];
  assign T427 = T126[5'h1d:5'h1d];
  assign T428 = T126[5'h1e:5'h1e];
  assign T429 = T126[5'h1f:5'h1f];
  assign T127 = T121 << 4'h9;
  assign T128 = T129 == 8'h0;
  assign T129 = load_wb_data[5'h1e:5'h17];
  assign T130 = T137 | T430;
  assign T430 = {2'h0, T131};
  assign T131 = T132 << 3'h6;
  assign T132 = T135 & T133;
  assign T133 = T134 ^ 1'h1;
  assign T134 = T121 == 23'h0;
  assign T135 = T136 == 2'h3;
  assign T136 = T137[4'h8:3'h7];
  assign T137 = T144 + T431;
  assign T431 = {1'h0, T138};
  assign T138 = T143 ? 8'h0 : T139;
  assign T139 = 8'h80 | T432;
  assign T432 = {6'h0, T140};
  assign T140 = T141 ? 2'h2 : 2'h1;
  assign T141 = T128 & T142;
  assign T142 = T134 ^ 1'h1;
  assign T143 = T128 & T134;
  assign T144 = T128 ? T145 : T433;
  assign T433 = {1'h0, T129};
  assign T145 = T134 ? 9'h0 : T146;
  assign T146 = {4'hf, T147};
  assign T147 = ~ T124;
  assign T148 = load_wb_data[5'h1f:5'h1f];
  assign T149 = io_dpath_dmem_resp_val ? T150 : load_wb_single;
  assign T150 = T152 | T151;
  assign T151 = T434 == 4'h6;
  assign T434 = {1'h0, io_dpath_dmem_resp_type};
  assign T152 = T435 == 4'h2;
  assign T435 = {1'h0, io_dpath_dmem_resp_type};
  assign T153 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_tag : load_wb_tag;
  assign T154 = T159 ? T158 : T155;
  assign T155 = T157 ? T156 : ex_ra3;
  assign T156 = io_dpath_inst[5'h1f:5'h1b];
  assign T157 = io_ctrl_valid & fp_decoder_io_sigs_ren3;
  assign T158 = io_dpath_inst[5'h18:5'h14];
  assign T159 = T162 & T160;
  assign T160 = T161 & fp_decoder_io_sigs_swap23;
  assign T161 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign T162 = io_ctrl_valid & fp_decoder_io_sigs_ren2;
  assign req_in2 = ex_rs2;
  assign ex_rs2 = regfile[ex_ra2];
  assign T163 = T165 ? T164 : ex_ra2;
  assign T164 = io_dpath_inst[5'h18:5'h14];
  assign T165 = T162 & T166;
  assign T166 = T168 & T167;
  assign T167 = fp_decoder_io_sigs_swap23 ^ 1'h1;
  assign T168 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign req_in1 = ex_rs1;
  assign ex_rs1 = regfile[ex_ra1];
  assign T169 = T174 ? T173 : T170;
  assign T170 = T172 ? T171 : ex_ra1;
  assign T171 = io_dpath_inst[5'h13:4'hf];
  assign T172 = io_ctrl_valid & fp_decoder_io_sigs_ren1;
  assign T173 = io_dpath_inst[5'h18:5'h14];
  assign T174 = T162 & fp_decoder_io_sigs_ldst;
  assign req_typ = T175;
  assign T175 = ex_reg_inst[5'h15:5'h14];
  assign req_rm = ex_rm;
  assign ex_rm = T177 ? io_dpath_fcsr_rm : T176;
  assign T176 = ex_reg_inst[4'he:4'hc];
  assign T177 = T178 == 3'h7;
  assign T178 = ex_reg_inst[4'he:4'hc];
  assign req_round = ex_ctrl_round;
  assign T179 = io_ctrl_valid ? fp_decoder_io_sigs_round : ex_ctrl_round;
  assign req_fma = ex_ctrl_fma;
  assign req_fastpipe = ex_ctrl_fastpipe;
  assign req_toint = ex_ctrl_toint;
  assign T180 = io_ctrl_valid ? fp_decoder_io_sigs_toint : ex_ctrl_toint;
  assign req_fromint = ex_ctrl_fromint;
  assign req_single = ex_ctrl_single;
  assign req_swap23 = ex_ctrl_swap23;
  assign T181 = io_ctrl_valid ? fp_decoder_io_sigs_swap23 : ex_ctrl_swap23;
  assign req_ren3 = ex_ctrl_ren3;
  assign T182 = io_ctrl_valid ? fp_decoder_io_sigs_ren3 : ex_ctrl_ren3;
  assign req_ren2 = ex_ctrl_ren2;
  assign T183 = io_ctrl_valid ? fp_decoder_io_sigs_ren2 : ex_ctrl_ren2;
  assign req_ren1 = ex_ctrl_ren1;
  assign T184 = io_ctrl_valid ? fp_decoder_io_sigs_ren1 : ex_ctrl_ren1;
  assign req_wen = ex_ctrl_wen;
  assign T185 = io_ctrl_valid ? fp_decoder_io_sigs_wen : ex_ctrl_wen;
  assign req_ldst = ex_ctrl_ldst;
  assign T186 = io_ctrl_valid ? fp_decoder_io_sigs_ldst : ex_ctrl_ldst;
  assign req_cmd = ex_ctrl_cmd;
  assign T187 = io_ctrl_valid ? fp_decoder_io_sigs_cmd : ex_ctrl_cmd;
  assign T188 = ex_reg_valid & ex_ctrl_fastpipe;
  assign T436 = {1'h0, io_dpath_fromint_data};
  assign T189 = ex_reg_valid & ex_ctrl_fromint;
  assign T190 = ex_reg_valid & T191;
  assign T191 = ex_ctrl_toint | T192;
  assign T192 = T193 == 5'h5;
  assign T193 = ex_ctrl_cmd & 5'hd;
  assign T194 = T196 & T195;
  assign T195 = ex_ctrl_single ^ 1'h1;
  assign T196 = ex_reg_valid & ex_ctrl_fma;
  assign T197 = T198 & ex_ctrl_single;
  assign T198 = ex_reg_valid & ex_ctrl_fma;
  assign io_dpath_toint_data = fpiu_io_out_bits_toint;
  assign io_dpath_store_data = fpiu_io_out_bits_store;
  assign io_dpath_fcsr_flags_bits = T199;
  assign T199 = T208 | T200;
  assign T200 = T207 ? wexc : 5'h0;
  assign wexc = T206 ? T204 : T201;
  assign T201 = T202 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc;
  assign T202 = T203[1'h0:1'h0];
  assign T203 = wsrc;
  assign T204 = T205 ? dfma_io_out_bits_exc : sfma_io_out_bits_exc;
  assign T205 = T203[1'h0:1'h0];
  assign T206 = T203[1'h1:1'h1];
  assign T207 = wen[1'h0:1'h0];
  assign T208 = wb_toint_valid ? wb_toint_exc : 5'h0;
  assign T209 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign T210 = ex_reg_valid ? ex_ctrl_toint : mem_ctrl_toint;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign T211 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign T437 = reset ? 1'h0 : T212;
  assign T212 = mem_reg_valid & T213;
  assign T213 = killm ^ 1'h1;
  assign io_dpath_fcsr_flags_valid = T214;
  assign T214 = wb_toint_valid | T215;
  assign T215 = wen[1'h0:1'h0];
  assign io_ctrl_sboard_clra = waddr;
  assign io_ctrl_sboard_clr = 1'h0;
  assign io_ctrl_sboard_set = T216;
  assign T216 = wb_reg_valid & R217;
  assign io_ctrl_dec_round = fp_decoder_io_sigs_round;
  assign io_ctrl_dec_fma = fp_decoder_io_sigs_fma;
  assign io_ctrl_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_ctrl_dec_toint = fp_decoder_io_sigs_toint;
  assign io_ctrl_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_ctrl_dec_single = fp_decoder_io_sigs_single;
  assign io_ctrl_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_ctrl_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_ctrl_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_ctrl_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_ctrl_dec_wen = fp_decoder_io_sigs_wen;
  assign io_ctrl_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_ctrl_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_ctrl_illegal_rm = T218;
  assign T218 = T219 & ex_ctrl_round;
  assign T219 = ex_rm[2'h2:2'h2];
  assign io_ctrl_nack_mem = write_port_busy;
  assign io_ctrl_fcsr_rdy = T220;
  assign T220 = fp_inflight ^ 1'h1;
  assign fp_inflight = T222 | T221;
  assign T221 = wen != 2'h0;
  assign T222 = wb_reg_valid & wb_ctrl_toint;
  FPUDecoder fp_decoder(
       .io_inst( io_dpath_inst ),
       .io_sigs_cmd( fp_decoder_io_sigs_cmd ),
       .io_sigs_ldst( fp_decoder_io_sigs_ldst ),
       .io_sigs_wen( fp_decoder_io_sigs_wen ),
       .io_sigs_ren1( fp_decoder_io_sigs_ren1 ),
       .io_sigs_ren2( fp_decoder_io_sigs_ren2 ),
       .io_sigs_ren3( fp_decoder_io_sigs_ren3 ),
       .io_sigs_swap23( fp_decoder_io_sigs_swap23 ),
       .io_sigs_single( fp_decoder_io_sigs_single ),
       .io_sigs_fromint( fp_decoder_io_sigs_fromint ),
       .io_sigs_toint( fp_decoder_io_sigs_toint ),
       .io_sigs_fastpipe( fp_decoder_io_sigs_fastpipe ),
       .io_sigs_fma( fp_decoder_io_sigs_fma ),
       .io_sigs_round( fp_decoder_io_sigs_round )
  );
  FPUFMAPipe_0 sfma(.clk(clk), .reset(reset),
       .io_in_valid( T197 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( sfma_io_out_bits_data ),
       .io_out_bits_exc( sfma_io_out_bits_exc )
  );
  FPUFMAPipe_1 dfma(.clk(clk), .reset(reset),
       .io_in_valid( T194 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( dfma_io_out_bits_data ),
       .io_out_bits_exc( dfma_io_out_bits_exc )
  );
  FPToInt fpiu(.clk(clk),
       .io_in_valid( T190 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_lt( fpiu_io_out_bits_lt ),
       .io_out_bits_store( fpiu_io_out_bits_store ),
       .io_out_bits_toint( fpiu_io_out_bits_toint ),
       .io_out_bits_exc( fpiu_io_out_bits_exc )
  );
  IntToFP ifpu(.clk(clk), .reset(reset),
       .io_in_valid( T189 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( T436 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( ifpu_io_out_bits_data ),
       .io_out_bits_exc( ifpu_io_out_bits_exc )
  );
  FPToFP fpmu(.clk(clk), .reset(reset),
       .io_in_valid( T188 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( fpmu_io_out_bits_data ),
       .io_out_bits_exc( fpmu_io_out_bits_exc ),
       .io_lt( fpiu_io_out_bits_lt )
  );

  always @(posedge clk) begin
    if (T83)
      regfile[T84] <= T223;
    if(T75) begin
      winfo_0 <= mem_winfo;
    end else if(T63) begin
      winfo_0 <= winfo_1;
    end
    if(T7) begin
      winfo_1 <= mem_winfo;
    end
    if(ex_reg_valid) begin
      mem_ctrl_single <= ex_ctrl_single;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_single <= fp_decoder_io_sigs_single;
    end
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_ctrl_valid;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fma <= ex_ctrl_fma;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fromint <= ex_ctrl_fromint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_ctrl_fastpipe;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if(ex_reg_valid) begin
      write_port_busy <= T27;
    end
    if(reset) begin
      wen <= 2'h0;
    end else if(T44) begin
      wen <= T42;
    end else begin
      wen <= T232;
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T61;
    end
    if(ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(io_ctrl_valid) begin
      ex_reg_inst <= io_dpath_inst;
    end
    if (load_wb)
      regfile[load_wb_tag] <= load_wb_data_recoded;
    if(io_dpath_dmem_resp_val) begin
      load_wb_data <= io_dpath_dmem_resp_data;
    end
    if(io_dpath_dmem_resp_val) begin
      load_wb_single <= T150;
    end
    load_wb <= io_dpath_dmem_resp_val;
    if(io_dpath_dmem_resp_val) begin
      load_wb_tag <= io_dpath_dmem_resp_tag;
    end
    if(T159) begin
      ex_ra3 <= T158;
    end else if(T157) begin
      ex_ra3 <= T156;
    end
    if(T165) begin
      ex_ra2 <= T164;
    end
    if(T174) begin
      ex_ra1 <= T173;
    end else if(T172) begin
      ex_ra1 <= T171;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_round <= fp_decoder_io_sigs_round;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren1 <= fp_decoder_io_sigs_ren1;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_wen <= fp_decoder_io_sigs_wen;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ldst <= fp_decoder_io_sigs_ldst;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_cmd <= fp_decoder_io_sigs_cmd;
    end
    if(mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if(ex_reg_valid) begin
      mem_ctrl_toint <= ex_ctrl_toint;
    end
    if(mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T212;
    end
    R217 <= 1'h0;
  end
endmodule

module Core(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[43:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [42:0] io_imem_btb_resp_bits_target,
    input [5:0] io_imem_btb_resp_bits_entry,
    input [6:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    //output io_imem_btb_update_bits_taken
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    output[42:0] io_imem_btb_update_bits_br_pc,
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output[42:0] io_imem_bht_update_bits_prediction_bits_target,
    output[5:0] io_imem_bht_update_bits_prediction_bits_entry,
    output[6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_bht_update_bits_pc,
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    output[42:0] io_imem_ras_update_bits_returnAddr,
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output[42:0] io_imem_ras_update_bits_prediction_bits_target,
    output[5:0] io_imem_ras_update_bits_prediction_bits_entry,
    output[6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[3:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output[43:0] io_dmem_req_bits_addr,
    output[7:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [3:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [3:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[3:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_imem_acquire_bits_payload_data,
    input  io_rocc_imem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_imem_acquire_bits_payload_subblock,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[135:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_manager_xact_id
    //output io_rocc_imem_grant_bits_payload_uncached
    //output[1:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_manager_xact_id,
    //output io_rocc_dmem_acquire_ready
    input  io_rocc_dmem_acquire_valid,
    input [1:0] io_rocc_dmem_acquire_bits_header_src,
    input [1:0] io_rocc_dmem_acquire_bits_header_dst,
    input [25:0] io_rocc_dmem_acquire_bits_payload_addr,
    input [1:0] io_rocc_dmem_acquire_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_acquire_bits_payload_data,
    input  io_rocc_dmem_acquire_bits_payload_uncached,
    input [1:0] io_rocc_dmem_acquire_bits_payload_a_type,
    input [128:0] io_rocc_dmem_acquire_bits_payload_subblock,
    input  io_rocc_dmem_grant_ready,
    //output io_rocc_dmem_grant_valid
    //output[1:0] io_rocc_dmem_grant_bits_header_src
    //output[1:0] io_rocc_dmem_grant_bits_header_dst
    //output[135:0] io_rocc_dmem_grant_bits_payload_data
    //output[1:0] io_rocc_dmem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_dmem_grant_bits_payload_manager_xact_id
    //output io_rocc_dmem_grant_bits_payload_uncached
    //output[1:0] io_rocc_dmem_grant_bits_payload_g_type
    //output io_rocc_dmem_finish_ready
    input  io_rocc_dmem_finish_valid,
    input [1:0] io_rocc_dmem_finish_bits_header_src,
    input [1:0] io_rocc_dmem_finish_bits_header_dst,
    input [3:0] io_rocc_dmem_finish_bits_payload_manager_xact_id,
    input  io_rocc_dmem_probe_ready,
    //output io_rocc_dmem_probe_valid
    //output[1:0] io_rocc_dmem_probe_bits_header_src
    //output[1:0] io_rocc_dmem_probe_bits_header_dst
    //output[25:0] io_rocc_dmem_probe_bits_payload_addr
    //output[1:0] io_rocc_dmem_probe_bits_payload_p_type
    //output io_rocc_dmem_release_ready
    input  io_rocc_dmem_release_valid,
    input [1:0] io_rocc_dmem_release_bits_header_src,
    input [1:0] io_rocc_dmem_release_bits_header_dst,
    input [25:0] io_rocc_dmem_release_bits_payload_addr,
    input [1:0] io_rocc_dmem_release_bits_payload_client_xact_id,
    input [135:0] io_rocc_dmem_release_bits_payload_data,
    input [2:0] io_rocc_dmem_release_bits_payload_r_type,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire[2:0] ctrl_io_dpath_sel_pc;
  wire ctrl_io_dpath_killd;
  wire ctrl_io_dpath_killm;
  wire ctrl_io_dpath_ren_1;
  wire ctrl_io_dpath_ren_0;
  wire ctrl_io_dpath_ex_ctrl_legal;
  wire ctrl_io_dpath_ex_ctrl_fp;
  wire ctrl_io_dpath_ex_ctrl_rocc;
  wire ctrl_io_dpath_ex_ctrl_branch;
  wire ctrl_io_dpath_ex_ctrl_jal;
  wire ctrl_io_dpath_ex_ctrl_jalr;
  wire ctrl_io_dpath_ex_ctrl_rxs2;
  wire ctrl_io_dpath_ex_ctrl_rxs1;
  wire[1:0] ctrl_io_dpath_ex_ctrl_sel_alu2;
  wire[1:0] ctrl_io_dpath_ex_ctrl_sel_alu1;
  wire[2:0] ctrl_io_dpath_ex_ctrl_sel_imm;
  wire ctrl_io_dpath_ex_ctrl_alu_dw;
  wire[3:0] ctrl_io_dpath_ex_ctrl_alu_fn;
  wire ctrl_io_dpath_ex_ctrl_mem;
  wire[4:0] ctrl_io_dpath_ex_ctrl_mem_cmd;
  wire[3:0] ctrl_io_dpath_ex_ctrl_mem_type;
  wire ctrl_io_dpath_ex_ctrl_rfs1;
  wire ctrl_io_dpath_ex_ctrl_rfs2;
  wire ctrl_io_dpath_ex_ctrl_rfs3;
  wire ctrl_io_dpath_ex_ctrl_wfd;
  wire ctrl_io_dpath_ex_ctrl_div;
  wire ctrl_io_dpath_ex_ctrl_wxd;
  wire[1:0] ctrl_io_dpath_ex_ctrl_csr;
  wire ctrl_io_dpath_ex_ctrl_fence_i;
  wire ctrl_io_dpath_ex_ctrl_sret;
  wire ctrl_io_dpath_ex_ctrl_scall;
  wire ctrl_io_dpath_ex_ctrl_fence;
  wire ctrl_io_dpath_ex_ctrl_amo;
  wire ctrl_io_dpath_mem_ctrl_legal;
  wire ctrl_io_dpath_mem_ctrl_fp;
  wire ctrl_io_dpath_mem_ctrl_rocc;
  wire ctrl_io_dpath_mem_ctrl_branch;
  wire ctrl_io_dpath_mem_ctrl_jal;
  wire ctrl_io_dpath_mem_ctrl_jalr;
  wire ctrl_io_dpath_mem_ctrl_rxs2;
  wire ctrl_io_dpath_mem_ctrl_rxs1;
  wire[1:0] ctrl_io_dpath_mem_ctrl_sel_alu2;
  wire[1:0] ctrl_io_dpath_mem_ctrl_sel_alu1;
  wire[2:0] ctrl_io_dpath_mem_ctrl_sel_imm;
  wire ctrl_io_dpath_mem_ctrl_alu_dw;
  wire[3:0] ctrl_io_dpath_mem_ctrl_alu_fn;
  wire ctrl_io_dpath_mem_ctrl_mem;
  wire[4:0] ctrl_io_dpath_mem_ctrl_mem_cmd;
  wire[3:0] ctrl_io_dpath_mem_ctrl_mem_type;
  wire ctrl_io_dpath_mem_ctrl_rfs1;
  wire ctrl_io_dpath_mem_ctrl_rfs2;
  wire ctrl_io_dpath_mem_ctrl_rfs3;
  wire ctrl_io_dpath_mem_ctrl_wfd;
  wire ctrl_io_dpath_mem_ctrl_div;
  wire ctrl_io_dpath_mem_ctrl_wxd;
  wire[1:0] ctrl_io_dpath_mem_ctrl_csr;
  wire ctrl_io_dpath_mem_ctrl_fence_i;
  wire ctrl_io_dpath_mem_ctrl_sret;
  wire ctrl_io_dpath_mem_ctrl_scall;
  wire ctrl_io_dpath_mem_ctrl_fence;
  wire ctrl_io_dpath_mem_ctrl_amo;
  wire[2:0] ctrl_io_dpath_csr;
  wire ctrl_io_dpath_sret;
  wire ctrl_io_dpath_ex_valid;
  wire ctrl_io_dpath_wb_wen;
  wire ctrl_io_dpath_bypass_1;
  wire ctrl_io_dpath_bypass_0;
  wire[1:0] ctrl_io_dpath_bypass_src_1;
  wire[1:0] ctrl_io_dpath_bypass_src_0;
  wire ctrl_io_dpath_ll_ready;
  wire ctrl_io_dpath_retire;
  wire ctrl_io_dpath_exception;
  wire[63:0] ctrl_io_dpath_cause;
  wire ctrl_io_dpath_badvaddr_wen;
  wire ctrl_io_imem_req_valid;
  wire ctrl_io_imem_resp_ready;
  wire ctrl_io_imem_btb_update_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_mask;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_bridx;
  wire[42:0] ctrl_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire ctrl_io_imem_btb_update_bits_isJump;
  wire ctrl_io_imem_btb_update_bits_isReturn;
  wire ctrl_io_imem_bht_update_valid;
  wire ctrl_io_imem_bht_update_bits_prediction_valid;
  wire ctrl_io_imem_bht_update_bits_prediction_bits_taken;
  wire ctrl_io_imem_bht_update_bits_prediction_bits_mask;
  wire ctrl_io_imem_bht_update_bits_prediction_bits_bridx;
  wire[42:0] ctrl_io_imem_bht_update_bits_prediction_bits_target;
  wire[5:0] ctrl_io_imem_bht_update_bits_prediction_bits_entry;
  wire[6:0] ctrl_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire[1:0] ctrl_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire ctrl_io_imem_bht_update_bits_taken;
  wire ctrl_io_imem_bht_update_bits_mispredict;
  wire ctrl_io_imem_ras_update_valid;
  wire ctrl_io_imem_ras_update_bits_isCall;
  wire ctrl_io_imem_ras_update_bits_isReturn;
  wire ctrl_io_imem_ras_update_bits_prediction_valid;
  wire ctrl_io_imem_ras_update_bits_prediction_bits_taken;
  wire ctrl_io_imem_ras_update_bits_prediction_bits_mask;
  wire ctrl_io_imem_ras_update_bits_prediction_bits_bridx;
  wire[42:0] ctrl_io_imem_ras_update_bits_prediction_bits_target;
  wire[5:0] ctrl_io_imem_ras_update_bits_prediction_bits_entry;
  wire[6:0] ctrl_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire[1:0] ctrl_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire ctrl_io_imem_invalidate;
  wire ctrl_io_dmem_req_valid;
  wire ctrl_io_dmem_req_bits_kill;
  wire[3:0] ctrl_io_dmem_req_bits_typ;
  wire ctrl_io_dmem_req_bits_phys;
  wire[4:0] ctrl_io_dmem_req_bits_cmd;
  wire ctrl_io_fpu_valid;
  wire ctrl_io_fpu_killx;
  wire ctrl_io_fpu_killm;
  wire ctrl_io_rocc_cmd_valid;
  wire ctrl_io_rocc_s;
  wire ctrl_io_rocc_exception;
  wire dpath_io_host_pcr_req_ready;
  wire dpath_io_host_pcr_rep_valid;
  wire[63:0] dpath_io_host_pcr_rep_bits;
  wire dpath_io_host_ipi_req_valid;
  wire dpath_io_host_ipi_req_bits;
  wire dpath_io_host_ipi_rep_ready;
  wire dpath_io_host_debug_stats_pcr;
  wire[31:0] dpath_io_ctrl_inst;
  wire dpath_io_ctrl_mem_br_taken;
  wire dpath_io_ctrl_mem_misprediction;
  wire dpath_io_ctrl_div_mul_rdy;
  wire dpath_io_ctrl_ll_wen;
  wire[4:0] dpath_io_ctrl_ll_waddr;
  wire[4:0] dpath_io_ctrl_ex_waddr;
  wire dpath_io_ctrl_mem_rs1_ra;
  wire[4:0] dpath_io_ctrl_mem_waddr;
  wire[4:0] dpath_io_ctrl_wb_waddr;
  wire[7:0] dpath_io_ctrl_status_ip;
  wire[7:0] dpath_io_ctrl_status_im;
  wire[6:0] dpath_io_ctrl_status_zero;
  wire dpath_io_ctrl_status_er;
  wire dpath_io_ctrl_status_vm;
  wire dpath_io_ctrl_status_s64;
  wire dpath_io_ctrl_status_u64;
  wire dpath_io_ctrl_status_ef;
  wire dpath_io_ctrl_status_pei;
  wire dpath_io_ctrl_status_ei;
  wire dpath_io_ctrl_status_ps;
  wire dpath_io_ctrl_status_s;
  wire dpath_io_ctrl_fp_sboard_clr;
  wire[4:0] dpath_io_ctrl_fp_sboard_clra;
  wire dpath_io_ctrl_csr_replay;
  wire[43:0] dpath_io_dmem_req_bits_addr;
  wire[7:0] dpath_io_dmem_req_bits_tag;
  wire[63:0] dpath_io_dmem_req_bits_data;
  wire[31:0] dpath_io_ptw_ptbr;
  wire dpath_io_ptw_invalidate;
  wire dpath_io_ptw_sret;
  wire[7:0] dpath_io_ptw_status_ip;
  wire[7:0] dpath_io_ptw_status_im;
  wire[6:0] dpath_io_ptw_status_zero;
  wire dpath_io_ptw_status_er;
  wire dpath_io_ptw_status_vm;
  wire dpath_io_ptw_status_s64;
  wire dpath_io_ptw_status_u64;
  wire dpath_io_ptw_status_ef;
  wire dpath_io_ptw_status_pei;
  wire dpath_io_ptw_status_ei;
  wire dpath_io_ptw_status_ps;
  wire dpath_io_ptw_status_s;
  wire[43:0] dpath_io_imem_req_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_target;
  wire[42:0] dpath_io_imem_btb_update_bits_br_pc;
  wire[42:0] dpath_io_imem_bht_update_bits_pc;
  wire[42:0] dpath_io_imem_ras_update_bits_returnAddr;
  wire[31:0] dpath_io_fpu_inst;
  wire[63:0] dpath_io_fpu_fromint_data;
  wire[2:0] dpath_io_fpu_fcsr_rm;
  wire dpath_io_fpu_dmem_resp_val;
  wire[2:0] dpath_io_fpu_dmem_resp_type;
  wire[4:0] dpath_io_fpu_dmem_resp_tag;
  wire[63:0] dpath_io_fpu_dmem_resp_data;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_funct;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs1;
  wire dpath_io_rocc_cmd_bits_inst_xd;
  wire dpath_io_rocc_cmd_bits_inst_xs1;
  wire dpath_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rd;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] dpath_io_rocc_cmd_bits_rs1;
  wire[63:0] dpath_io_rocc_cmd_bits_rs2;
  wire FPU_io_ctrl_fcsr_rdy;
  wire FPU_io_ctrl_nack_mem;
  wire FPU_io_ctrl_illegal_rm;
  wire[4:0] FPU_io_ctrl_dec_cmd;
  wire FPU_io_ctrl_dec_ldst;
  wire FPU_io_ctrl_dec_wen;
  wire FPU_io_ctrl_dec_ren1;
  wire FPU_io_ctrl_dec_ren2;
  wire FPU_io_ctrl_dec_ren3;
  wire FPU_io_ctrl_dec_swap23;
  wire FPU_io_ctrl_dec_single;
  wire FPU_io_ctrl_dec_fromint;
  wire FPU_io_ctrl_dec_toint;
  wire FPU_io_ctrl_dec_fastpipe;
  wire FPU_io_ctrl_dec_fma;
  wire FPU_io_ctrl_dec_round;
  wire FPU_io_ctrl_sboard_set;
  wire FPU_io_ctrl_sboard_clr;
  wire[4:0] FPU_io_ctrl_sboard_clra;
  wire FPU_io_dpath_fcsr_flags_valid;
  wire[4:0] FPU_io_dpath_fcsr_flags_bits;
  wire[63:0] FPU_io_dpath_store_data;
  wire[63:0] FPU_io_dpath_toint_data;


  assign io_rocc_exception = ctrl_io_rocc_exception;
//  assign io_rocc_pptw_sret = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_s = {1{$random}};
//  assign io_rocc_pptw_status_ps = {1{$random}};
//  assign io_rocc_pptw_status_ei = {1{$random}};
//  assign io_rocc_pptw_status_pei = {1{$random}};
//  assign io_rocc_pptw_status_ef = {1{$random}};
//  assign io_rocc_pptw_status_u64 = {1{$random}};
//  assign io_rocc_pptw_status_s64 = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_er = {1{$random}};
//  assign io_rocc_pptw_status_zero = {1{$random}};
//  assign io_rocc_pptw_status_im = {1{$random}};
//  assign io_rocc_pptw_status_ip = {1{$random}};
//  assign io_rocc_pptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_pptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_sret = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_s = {1{$random}};
//  assign io_rocc_dptw_status_ps = {1{$random}};
//  assign io_rocc_dptw_status_ei = {1{$random}};
//  assign io_rocc_dptw_status_pei = {1{$random}};
//  assign io_rocc_dptw_status_ef = {1{$random}};
//  assign io_rocc_dptw_status_u64 = {1{$random}};
//  assign io_rocc_dptw_status_s64 = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_er = {1{$random}};
//  assign io_rocc_dptw_status_zero = {1{$random}};
//  assign io_rocc_dptw_status_im = {1{$random}};
//  assign io_rocc_dptw_status_ip = {1{$random}};
//  assign io_rocc_dptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_dptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_sret = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_s = {1{$random}};
//  assign io_rocc_iptw_status_ps = {1{$random}};
//  assign io_rocc_iptw_status_ei = {1{$random}};
//  assign io_rocc_iptw_status_pei = {1{$random}};
//  assign io_rocc_iptw_status_ef = {1{$random}};
//  assign io_rocc_iptw_status_u64 = {1{$random}};
//  assign io_rocc_iptw_status_s64 = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_er = {1{$random}};
//  assign io_rocc_iptw_status_zero = {1{$random}};
//  assign io_rocc_iptw_status_im = {1{$random}};
//  assign io_rocc_iptw_status_ip = {1{$random}};
//  assign io_rocc_iptw_resp_bits_perm = {1{$random}};
//  assign io_rocc_iptw_resp_bits_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_release_ready = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_p_type = {1{$random}};
//  assign io_rocc_dmem_probe_bits_payload_addr = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_probe_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_probe_valid = {1{$random}};
//  assign io_rocc_dmem_finish_ready = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_dmem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_dmem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_dmem_grant_valid = {1{$random}};
//  assign io_rocc_dmem_acquire_ready = {1{$random}};
//  assign io_rocc_imem_finish_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_uncached = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_payload_data = {5{$random}};
//  assign io_rocc_imem_grant_bits_header_dst = {1{$random}};
//  assign io_rocc_imem_grant_bits_header_src = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
  assign io_rocc_s = ctrl_io_rocc_s;
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_ptw_req_bits = {1{$random}};
//  assign io_rocc_mem_ptw_req_valid = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_data_subword = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
  assign io_rocc_cmd_bits_rs2 = dpath_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = dpath_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = dpath_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = dpath_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = dpath_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = dpath_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = dpath_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = dpath_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = dpath_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = dpath_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = ctrl_io_rocc_cmd_valid;
  assign io_ptw_status_s = dpath_io_ptw_status_s;
  assign io_ptw_status_ps = dpath_io_ptw_status_ps;
  assign io_ptw_status_ei = dpath_io_ptw_status_ei;
  assign io_ptw_status_pei = dpath_io_ptw_status_pei;
  assign io_ptw_status_ef = dpath_io_ptw_status_ef;
  assign io_ptw_status_u64 = dpath_io_ptw_status_u64;
  assign io_ptw_status_s64 = dpath_io_ptw_status_s64;
  assign io_ptw_status_vm = dpath_io_ptw_status_vm;
  assign io_ptw_status_er = dpath_io_ptw_status_er;
  assign io_ptw_status_zero = dpath_io_ptw_status_zero;
  assign io_ptw_status_im = dpath_io_ptw_status_im;
  assign io_ptw_status_ip = dpath_io_ptw_status_ip;
  assign io_ptw_sret = dpath_io_ptw_sret;
  assign io_ptw_invalidate = dpath_io_ptw_invalidate;
  assign io_ptw_ptbr = dpath_io_ptw_ptbr;
//  assign io_dmem_ptw_sret = {1{$random}};
//  assign io_dmem_ptw_invalidate = {1{$random}};
//  assign io_dmem_ptw_status_s = {1{$random}};
//  assign io_dmem_ptw_status_ps = {1{$random}};
//  assign io_dmem_ptw_status_ei = {1{$random}};
//  assign io_dmem_ptw_status_pei = {1{$random}};
//  assign io_dmem_ptw_status_ef = {1{$random}};
//  assign io_dmem_ptw_status_u64 = {1{$random}};
//  assign io_dmem_ptw_status_s64 = {1{$random}};
//  assign io_dmem_ptw_status_vm = {1{$random}};
//  assign io_dmem_ptw_status_er = {1{$random}};
//  assign io_dmem_ptw_status_zero = {1{$random}};
//  assign io_dmem_ptw_status_im = {1{$random}};
//  assign io_dmem_ptw_status_ip = {1{$random}};
//  assign io_dmem_ptw_resp_bits_perm = {1{$random}};
//  assign io_dmem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_dmem_ptw_resp_bits_error = {1{$random}};
//  assign io_dmem_ptw_resp_valid = {1{$random}};
//  assign io_dmem_ptw_req_ready = {1{$random}};
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_cmd = ctrl_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_tag = dpath_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_phys = ctrl_io_dmem_req_bits_phys;
  assign io_dmem_req_bits_typ = ctrl_io_dmem_req_bits_typ;
  assign io_dmem_req_bits_kill = ctrl_io_dmem_req_bits_kill;
  assign io_dmem_req_valid = ctrl_io_dmem_req_valid;
  assign io_imem_invalidate = ctrl_io_imem_invalidate;
//  assign io_imem_ptw_sret = {1{$random}};
//  assign io_imem_ptw_invalidate = {1{$random}};
//  assign io_imem_ptw_status_s = {1{$random}};
//  assign io_imem_ptw_status_ps = {1{$random}};
//  assign io_imem_ptw_status_ei = {1{$random}};
//  assign io_imem_ptw_status_pei = {1{$random}};
//  assign io_imem_ptw_status_ef = {1{$random}};
//  assign io_imem_ptw_status_u64 = {1{$random}};
//  assign io_imem_ptw_status_s64 = {1{$random}};
//  assign io_imem_ptw_status_vm = {1{$random}};
//  assign io_imem_ptw_status_er = {1{$random}};
//  assign io_imem_ptw_status_zero = {1{$random}};
//  assign io_imem_ptw_status_im = {1{$random}};
//  assign io_imem_ptw_status_ip = {1{$random}};
//  assign io_imem_ptw_resp_bits_perm = {1{$random}};
//  assign io_imem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_imem_ptw_resp_bits_error = {1{$random}};
//  assign io_imem_ptw_resp_valid = {1{$random}};
//  assign io_imem_ptw_req_ready = {1{$random}};
  assign io_imem_ras_update_bits_prediction_bits_bht_value = ctrl_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = ctrl_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_entry = ctrl_io_imem_ras_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_target = ctrl_io_imem_ras_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_bridx = ctrl_io_imem_ras_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_mask = ctrl_io_imem_ras_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_taken = ctrl_io_imem_ras_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_valid = ctrl_io_imem_ras_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_returnAddr = dpath_io_imem_ras_update_bits_returnAddr;
  assign io_imem_ras_update_bits_isReturn = ctrl_io_imem_ras_update_bits_isReturn;
  assign io_imem_ras_update_bits_isCall = ctrl_io_imem_ras_update_bits_isCall;
  assign io_imem_ras_update_valid = ctrl_io_imem_ras_update_valid;
  assign io_imem_bht_update_bits_mispredict = ctrl_io_imem_bht_update_bits_mispredict;
  assign io_imem_bht_update_bits_taken = ctrl_io_imem_bht_update_bits_taken;
  assign io_imem_bht_update_bits_pc = dpath_io_imem_bht_update_bits_pc;
  assign io_imem_bht_update_bits_prediction_bits_bht_value = ctrl_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = ctrl_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_entry = ctrl_io_imem_bht_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_target = ctrl_io_imem_bht_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_bridx = ctrl_io_imem_bht_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_mask = ctrl_io_imem_bht_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_taken = ctrl_io_imem_bht_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_valid = ctrl_io_imem_bht_update_bits_prediction_valid;
  assign io_imem_bht_update_valid = ctrl_io_imem_bht_update_valid;
  assign io_imem_btb_update_bits_br_pc = dpath_io_imem_btb_update_bits_br_pc;
  assign io_imem_btb_update_bits_isReturn = ctrl_io_imem_btb_update_bits_isReturn;
  assign io_imem_btb_update_bits_isJump = ctrl_io_imem_btb_update_bits_isJump;
//  assign io_imem_btb_update_bits_taken = {1{$random}};
  assign io_imem_btb_update_bits_target = dpath_io_imem_btb_update_bits_target;
  assign io_imem_btb_update_bits_pc = dpath_io_imem_btb_update_bits_pc;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = ctrl_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = ctrl_io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_btb_update_bits_prediction_bits_bridx = ctrl_io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_btb_update_bits_prediction_bits_mask = ctrl_io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_btb_update_bits_prediction_bits_taken = ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_btb_update_bits_prediction_valid = ctrl_io_imem_btb_update_bits_prediction_valid;
  assign io_imem_btb_update_valid = ctrl_io_imem_btb_update_valid;
  assign io_imem_resp_ready = ctrl_io_imem_resp_ready;
  assign io_imem_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign io_imem_req_valid = ctrl_io_imem_req_valid;
  assign io_host_debug_stats_pcr = dpath_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = dpath_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = dpath_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = dpath_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = dpath_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = dpath_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = dpath_io_host_pcr_req_ready;
  Control ctrl(.clk(clk), .reset(reset),
       .io_dpath_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_dpath_killd( ctrl_io_dpath_killd ),
       .io_dpath_killm( ctrl_io_dpath_killm ),
       .io_dpath_ren_1( ctrl_io_dpath_ren_1 ),
       .io_dpath_ren_0( ctrl_io_dpath_ren_0 ),
       .io_dpath_ex_ctrl_legal( ctrl_io_dpath_ex_ctrl_legal ),
       .io_dpath_ex_ctrl_fp( ctrl_io_dpath_ex_ctrl_fp ),
       .io_dpath_ex_ctrl_rocc( ctrl_io_dpath_ex_ctrl_rocc ),
       .io_dpath_ex_ctrl_branch( ctrl_io_dpath_ex_ctrl_branch ),
       .io_dpath_ex_ctrl_jal( ctrl_io_dpath_ex_ctrl_jal ),
       .io_dpath_ex_ctrl_jalr( ctrl_io_dpath_ex_ctrl_jalr ),
       .io_dpath_ex_ctrl_rxs2( ctrl_io_dpath_ex_ctrl_rxs2 ),
       .io_dpath_ex_ctrl_rxs1( ctrl_io_dpath_ex_ctrl_rxs1 ),
       .io_dpath_ex_ctrl_sel_alu2( ctrl_io_dpath_ex_ctrl_sel_alu2 ),
       .io_dpath_ex_ctrl_sel_alu1( ctrl_io_dpath_ex_ctrl_sel_alu1 ),
       .io_dpath_ex_ctrl_sel_imm( ctrl_io_dpath_ex_ctrl_sel_imm ),
       .io_dpath_ex_ctrl_alu_dw( ctrl_io_dpath_ex_ctrl_alu_dw ),
       .io_dpath_ex_ctrl_alu_fn( ctrl_io_dpath_ex_ctrl_alu_fn ),
       .io_dpath_ex_ctrl_mem( ctrl_io_dpath_ex_ctrl_mem ),
       .io_dpath_ex_ctrl_mem_cmd( ctrl_io_dpath_ex_ctrl_mem_cmd ),
       .io_dpath_ex_ctrl_mem_type( ctrl_io_dpath_ex_ctrl_mem_type ),
       .io_dpath_ex_ctrl_rfs1( ctrl_io_dpath_ex_ctrl_rfs1 ),
       .io_dpath_ex_ctrl_rfs2( ctrl_io_dpath_ex_ctrl_rfs2 ),
       .io_dpath_ex_ctrl_rfs3( ctrl_io_dpath_ex_ctrl_rfs3 ),
       .io_dpath_ex_ctrl_wfd( ctrl_io_dpath_ex_ctrl_wfd ),
       .io_dpath_ex_ctrl_div( ctrl_io_dpath_ex_ctrl_div ),
       .io_dpath_ex_ctrl_wxd( ctrl_io_dpath_ex_ctrl_wxd ),
       .io_dpath_ex_ctrl_csr( ctrl_io_dpath_ex_ctrl_csr ),
       .io_dpath_ex_ctrl_fence_i( ctrl_io_dpath_ex_ctrl_fence_i ),
       .io_dpath_ex_ctrl_sret( ctrl_io_dpath_ex_ctrl_sret ),
       .io_dpath_ex_ctrl_scall( ctrl_io_dpath_ex_ctrl_scall ),
       .io_dpath_ex_ctrl_fence( ctrl_io_dpath_ex_ctrl_fence ),
       .io_dpath_ex_ctrl_amo( ctrl_io_dpath_ex_ctrl_amo ),
       .io_dpath_mem_ctrl_legal( ctrl_io_dpath_mem_ctrl_legal ),
       .io_dpath_mem_ctrl_fp( ctrl_io_dpath_mem_ctrl_fp ),
       .io_dpath_mem_ctrl_rocc( ctrl_io_dpath_mem_ctrl_rocc ),
       .io_dpath_mem_ctrl_branch( ctrl_io_dpath_mem_ctrl_branch ),
       .io_dpath_mem_ctrl_jal( ctrl_io_dpath_mem_ctrl_jal ),
       .io_dpath_mem_ctrl_jalr( ctrl_io_dpath_mem_ctrl_jalr ),
       .io_dpath_mem_ctrl_rxs2( ctrl_io_dpath_mem_ctrl_rxs2 ),
       .io_dpath_mem_ctrl_rxs1( ctrl_io_dpath_mem_ctrl_rxs1 ),
       .io_dpath_mem_ctrl_sel_alu2( ctrl_io_dpath_mem_ctrl_sel_alu2 ),
       .io_dpath_mem_ctrl_sel_alu1( ctrl_io_dpath_mem_ctrl_sel_alu1 ),
       .io_dpath_mem_ctrl_sel_imm( ctrl_io_dpath_mem_ctrl_sel_imm ),
       .io_dpath_mem_ctrl_alu_dw( ctrl_io_dpath_mem_ctrl_alu_dw ),
       .io_dpath_mem_ctrl_alu_fn( ctrl_io_dpath_mem_ctrl_alu_fn ),
       .io_dpath_mem_ctrl_mem( ctrl_io_dpath_mem_ctrl_mem ),
       .io_dpath_mem_ctrl_mem_cmd( ctrl_io_dpath_mem_ctrl_mem_cmd ),
       .io_dpath_mem_ctrl_mem_type( ctrl_io_dpath_mem_ctrl_mem_type ),
       .io_dpath_mem_ctrl_rfs1( ctrl_io_dpath_mem_ctrl_rfs1 ),
       .io_dpath_mem_ctrl_rfs2( ctrl_io_dpath_mem_ctrl_rfs2 ),
       .io_dpath_mem_ctrl_rfs3( ctrl_io_dpath_mem_ctrl_rfs3 ),
       .io_dpath_mem_ctrl_wfd( ctrl_io_dpath_mem_ctrl_wfd ),
       .io_dpath_mem_ctrl_div( ctrl_io_dpath_mem_ctrl_div ),
       .io_dpath_mem_ctrl_wxd( ctrl_io_dpath_mem_ctrl_wxd ),
       .io_dpath_mem_ctrl_csr( ctrl_io_dpath_mem_ctrl_csr ),
       .io_dpath_mem_ctrl_fence_i( ctrl_io_dpath_mem_ctrl_fence_i ),
       .io_dpath_mem_ctrl_sret( ctrl_io_dpath_mem_ctrl_sret ),
       .io_dpath_mem_ctrl_scall( ctrl_io_dpath_mem_ctrl_scall ),
       .io_dpath_mem_ctrl_fence( ctrl_io_dpath_mem_ctrl_fence ),
       .io_dpath_mem_ctrl_amo( ctrl_io_dpath_mem_ctrl_amo ),
       .io_dpath_csr( ctrl_io_dpath_csr ),
       .io_dpath_sret( ctrl_io_dpath_sret ),
       .io_dpath_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_dpath_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_dpath_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_dpath_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_dpath_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_dpath_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_dpath_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_dpath_retire( ctrl_io_dpath_retire ),
       .io_dpath_exception( ctrl_io_dpath_exception ),
       .io_dpath_cause( ctrl_io_dpath_cause ),
       .io_dpath_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_dpath_inst( dpath_io_ctrl_inst ),
       .io_dpath_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_dpath_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_dpath_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_dpath_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_dpath_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_dpath_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_dpath_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_dpath_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_dpath_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_dpath_status_ip( dpath_io_ctrl_status_ip ),
       .io_dpath_status_im( dpath_io_ctrl_status_im ),
       .io_dpath_status_zero( dpath_io_ctrl_status_zero ),
       .io_dpath_status_er( dpath_io_ctrl_status_er ),
       .io_dpath_status_vm( dpath_io_ctrl_status_vm ),
       .io_dpath_status_s64( dpath_io_ctrl_status_s64 ),
       .io_dpath_status_u64( dpath_io_ctrl_status_u64 ),
       .io_dpath_status_ef( dpath_io_ctrl_status_ef ),
       .io_dpath_status_pei( dpath_io_ctrl_status_pei ),
       .io_dpath_status_ei( dpath_io_ctrl_status_ei ),
       .io_dpath_status_ps( dpath_io_ctrl_status_ps ),
       .io_dpath_status_s( dpath_io_ctrl_status_s ),
       .io_dpath_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_dpath_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_dpath_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_imem_req_valid( ctrl_io_imem_req_valid ),
       //.io_imem_req_bits_pc(  )
       .io_imem_resp_ready( ctrl_io_imem_resp_ready ),
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data_0( io_imem_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( io_imem_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( io_imem_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( io_imem_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( io_imem_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( ctrl_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( ctrl_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( ctrl_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_mask( ctrl_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_imem_btb_update_bits_prediction_bits_bridx( ctrl_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_imem_btb_update_bits_prediction_bits_target( ctrl_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( ctrl_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( ctrl_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( ctrl_io_imem_btb_update_bits_prediction_bits_bht_value ),
       //.io_imem_btb_update_bits_pc(  )
       //.io_imem_btb_update_bits_target(  )
       //.io_imem_btb_update_bits_taken(  )
       .io_imem_btb_update_bits_isJump( ctrl_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isReturn( ctrl_io_imem_btb_update_bits_isReturn ),
       //.io_imem_btb_update_bits_br_pc(  )
       .io_imem_bht_update_valid( ctrl_io_imem_bht_update_valid ),
       .io_imem_bht_update_bits_prediction_valid( ctrl_io_imem_bht_update_bits_prediction_valid ),
       .io_imem_bht_update_bits_prediction_bits_taken( ctrl_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_imem_bht_update_bits_prediction_bits_mask( ctrl_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_imem_bht_update_bits_prediction_bits_bridx( ctrl_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_imem_bht_update_bits_prediction_bits_target( ctrl_io_imem_bht_update_bits_prediction_bits_target ),
       .io_imem_bht_update_bits_prediction_bits_entry( ctrl_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_imem_bht_update_bits_prediction_bits_bht_history( ctrl_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_imem_bht_update_bits_prediction_bits_bht_value( ctrl_io_imem_bht_update_bits_prediction_bits_bht_value ),
       //.io_imem_bht_update_bits_pc(  )
       .io_imem_bht_update_bits_taken( ctrl_io_imem_bht_update_bits_taken ),
       .io_imem_bht_update_bits_mispredict( ctrl_io_imem_bht_update_bits_mispredict ),
       .io_imem_ras_update_valid( ctrl_io_imem_ras_update_valid ),
       .io_imem_ras_update_bits_isCall( ctrl_io_imem_ras_update_bits_isCall ),
       .io_imem_ras_update_bits_isReturn( ctrl_io_imem_ras_update_bits_isReturn ),
       //.io_imem_ras_update_bits_returnAddr(  )
       .io_imem_ras_update_bits_prediction_valid( ctrl_io_imem_ras_update_bits_prediction_valid ),
       .io_imem_ras_update_bits_prediction_bits_taken( ctrl_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_imem_ras_update_bits_prediction_bits_mask( ctrl_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_imem_ras_update_bits_prediction_bits_bridx( ctrl_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_imem_ras_update_bits_prediction_bits_target( ctrl_io_imem_ras_update_bits_prediction_bits_target ),
       .io_imem_ras_update_bits_prediction_bits_entry( ctrl_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_imem_ras_update_bits_prediction_bits_bht_history( ctrl_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_imem_ras_update_bits_prediction_bits_bht_value( ctrl_io_imem_ras_update_bits_prediction_bits_bht_value ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( ctrl_io_imem_invalidate ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       .io_dmem_req_valid( ctrl_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( ctrl_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( ctrl_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( ctrl_io_dmem_req_bits_phys ),
       //.io_dmem_req_bits_addr(  )
       //.io_dmem_req_bits_tag(  )
       .io_dmem_req_bits_cmd( ctrl_io_dmem_req_bits_cmd ),
       //.io_dmem_req_bits_data(  )
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_fpu_valid( ctrl_io_fpu_valid ),
       .io_fpu_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_fpu_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_fpu_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_fpu_killx( ctrl_io_fpu_killx ),
       .io_fpu_killm( ctrl_io_fpu_killm ),
       .io_fpu_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_fpu_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_fpu_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_fpu_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_fpu_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_fpu_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_fpu_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_fpu_dec_single( FPU_io_ctrl_dec_single ),
       .io_fpu_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_fpu_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_fpu_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_fpu_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_fpu_dec_round( FPU_io_ctrl_dec_round ),
       .io_fpu_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_fpu_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_fpu_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( ctrl_io_rocc_cmd_valid ),
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( ctrl_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_manager_xact_id( io_rocc_imem_finish_bits_payload_manager_xact_id ),
       //.io_rocc_dmem_acquire_ready(  )
       .io_rocc_dmem_acquire_valid( io_rocc_dmem_acquire_valid ),
       .io_rocc_dmem_acquire_bits_header_src( io_rocc_dmem_acquire_bits_header_src ),
       .io_rocc_dmem_acquire_bits_header_dst( io_rocc_dmem_acquire_bits_header_dst ),
       .io_rocc_dmem_acquire_bits_payload_addr( io_rocc_dmem_acquire_bits_payload_addr ),
       .io_rocc_dmem_acquire_bits_payload_client_xact_id( io_rocc_dmem_acquire_bits_payload_client_xact_id ),
       .io_rocc_dmem_acquire_bits_payload_data( io_rocc_dmem_acquire_bits_payload_data ),
       .io_rocc_dmem_acquire_bits_payload_uncached( io_rocc_dmem_acquire_bits_payload_uncached ),
       .io_rocc_dmem_acquire_bits_payload_a_type( io_rocc_dmem_acquire_bits_payload_a_type ),
       .io_rocc_dmem_acquire_bits_payload_subblock( io_rocc_dmem_acquire_bits_payload_subblock ),
       .io_rocc_dmem_grant_ready( io_rocc_dmem_grant_ready ),
       //.io_rocc_dmem_grant_valid(  )
       //.io_rocc_dmem_grant_bits_header_src(  )
       //.io_rocc_dmem_grant_bits_header_dst(  )
       //.io_rocc_dmem_grant_bits_payload_data(  )
       //.io_rocc_dmem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_uncached(  )
       //.io_rocc_dmem_grant_bits_payload_g_type(  )
       //.io_rocc_dmem_finish_ready(  )
       .io_rocc_dmem_finish_valid( io_rocc_dmem_finish_valid ),
       .io_rocc_dmem_finish_bits_header_src( io_rocc_dmem_finish_bits_header_src ),
       .io_rocc_dmem_finish_bits_header_dst( io_rocc_dmem_finish_bits_header_dst ),
       .io_rocc_dmem_finish_bits_payload_manager_xact_id( io_rocc_dmem_finish_bits_payload_manager_xact_id ),
       .io_rocc_dmem_probe_ready( io_rocc_dmem_probe_ready ),
       //.io_rocc_dmem_probe_valid(  )
       //.io_rocc_dmem_probe_bits_header_src(  )
       //.io_rocc_dmem_probe_bits_header_dst(  )
       //.io_rocc_dmem_probe_bits_payload_addr(  )
       //.io_rocc_dmem_probe_bits_payload_p_type(  )
       //.io_rocc_dmem_release_ready(  )
       .io_rocc_dmem_release_valid( io_rocc_dmem_release_valid ),
       .io_rocc_dmem_release_bits_header_src( io_rocc_dmem_release_bits_header_src ),
       .io_rocc_dmem_release_bits_header_dst( io_rocc_dmem_release_bits_header_dst ),
       .io_rocc_dmem_release_bits_payload_addr( io_rocc_dmem_release_bits_payload_addr ),
       .io_rocc_dmem_release_bits_payload_client_xact_id( io_rocc_dmem_release_bits_payload_client_xact_id ),
       .io_rocc_dmem_release_bits_payload_data( io_rocc_dmem_release_bits_payload_data ),
       .io_rocc_dmem_release_bits_payload_r_type( io_rocc_dmem_release_bits_payload_r_type ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( ctrl_io_rocc_exception )
  );
  Datapath dpath(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( dpath_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( dpath_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( dpath_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( dpath_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( dpath_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( dpath_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( dpath_io_host_debug_stats_pcr ),
       .io_ctrl_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_ctrl_killd( ctrl_io_dpath_killd ),
       .io_ctrl_killm( ctrl_io_dpath_killm ),
       .io_ctrl_ren_1( ctrl_io_dpath_ren_1 ),
       .io_ctrl_ren_0( ctrl_io_dpath_ren_0 ),
       .io_ctrl_ex_ctrl_legal( ctrl_io_dpath_ex_ctrl_legal ),
       .io_ctrl_ex_ctrl_fp( ctrl_io_dpath_ex_ctrl_fp ),
       .io_ctrl_ex_ctrl_rocc( ctrl_io_dpath_ex_ctrl_rocc ),
       .io_ctrl_ex_ctrl_branch( ctrl_io_dpath_ex_ctrl_branch ),
       .io_ctrl_ex_ctrl_jal( ctrl_io_dpath_ex_ctrl_jal ),
       .io_ctrl_ex_ctrl_jalr( ctrl_io_dpath_ex_ctrl_jalr ),
       .io_ctrl_ex_ctrl_rxs2( ctrl_io_dpath_ex_ctrl_rxs2 ),
       .io_ctrl_ex_ctrl_rxs1( ctrl_io_dpath_ex_ctrl_rxs1 ),
       .io_ctrl_ex_ctrl_sel_alu2( ctrl_io_dpath_ex_ctrl_sel_alu2 ),
       .io_ctrl_ex_ctrl_sel_alu1( ctrl_io_dpath_ex_ctrl_sel_alu1 ),
       .io_ctrl_ex_ctrl_sel_imm( ctrl_io_dpath_ex_ctrl_sel_imm ),
       .io_ctrl_ex_ctrl_alu_dw( ctrl_io_dpath_ex_ctrl_alu_dw ),
       .io_ctrl_ex_ctrl_alu_fn( ctrl_io_dpath_ex_ctrl_alu_fn ),
       .io_ctrl_ex_ctrl_mem( ctrl_io_dpath_ex_ctrl_mem ),
       .io_ctrl_ex_ctrl_mem_cmd( ctrl_io_dpath_ex_ctrl_mem_cmd ),
       .io_ctrl_ex_ctrl_mem_type( ctrl_io_dpath_ex_ctrl_mem_type ),
       .io_ctrl_ex_ctrl_rfs1( ctrl_io_dpath_ex_ctrl_rfs1 ),
       .io_ctrl_ex_ctrl_rfs2( ctrl_io_dpath_ex_ctrl_rfs2 ),
       .io_ctrl_ex_ctrl_rfs3( ctrl_io_dpath_ex_ctrl_rfs3 ),
       .io_ctrl_ex_ctrl_wfd( ctrl_io_dpath_ex_ctrl_wfd ),
       .io_ctrl_ex_ctrl_div( ctrl_io_dpath_ex_ctrl_div ),
       .io_ctrl_ex_ctrl_wxd( ctrl_io_dpath_ex_ctrl_wxd ),
       .io_ctrl_ex_ctrl_csr( ctrl_io_dpath_ex_ctrl_csr ),
       .io_ctrl_ex_ctrl_fence_i( ctrl_io_dpath_ex_ctrl_fence_i ),
       .io_ctrl_ex_ctrl_sret( ctrl_io_dpath_ex_ctrl_sret ),
       .io_ctrl_ex_ctrl_scall( ctrl_io_dpath_ex_ctrl_scall ),
       .io_ctrl_ex_ctrl_fence( ctrl_io_dpath_ex_ctrl_fence ),
       .io_ctrl_ex_ctrl_amo( ctrl_io_dpath_ex_ctrl_amo ),
       .io_ctrl_mem_ctrl_legal( ctrl_io_dpath_mem_ctrl_legal ),
       .io_ctrl_mem_ctrl_fp( ctrl_io_dpath_mem_ctrl_fp ),
       .io_ctrl_mem_ctrl_rocc( ctrl_io_dpath_mem_ctrl_rocc ),
       .io_ctrl_mem_ctrl_branch( ctrl_io_dpath_mem_ctrl_branch ),
       .io_ctrl_mem_ctrl_jal( ctrl_io_dpath_mem_ctrl_jal ),
       .io_ctrl_mem_ctrl_jalr( ctrl_io_dpath_mem_ctrl_jalr ),
       .io_ctrl_mem_ctrl_rxs2( ctrl_io_dpath_mem_ctrl_rxs2 ),
       .io_ctrl_mem_ctrl_rxs1( ctrl_io_dpath_mem_ctrl_rxs1 ),
       .io_ctrl_mem_ctrl_sel_alu2( ctrl_io_dpath_mem_ctrl_sel_alu2 ),
       .io_ctrl_mem_ctrl_sel_alu1( ctrl_io_dpath_mem_ctrl_sel_alu1 ),
       .io_ctrl_mem_ctrl_sel_imm( ctrl_io_dpath_mem_ctrl_sel_imm ),
       .io_ctrl_mem_ctrl_alu_dw( ctrl_io_dpath_mem_ctrl_alu_dw ),
       .io_ctrl_mem_ctrl_alu_fn( ctrl_io_dpath_mem_ctrl_alu_fn ),
       .io_ctrl_mem_ctrl_mem( ctrl_io_dpath_mem_ctrl_mem ),
       .io_ctrl_mem_ctrl_mem_cmd( ctrl_io_dpath_mem_ctrl_mem_cmd ),
       .io_ctrl_mem_ctrl_mem_type( ctrl_io_dpath_mem_ctrl_mem_type ),
       .io_ctrl_mem_ctrl_rfs1( ctrl_io_dpath_mem_ctrl_rfs1 ),
       .io_ctrl_mem_ctrl_rfs2( ctrl_io_dpath_mem_ctrl_rfs2 ),
       .io_ctrl_mem_ctrl_rfs3( ctrl_io_dpath_mem_ctrl_rfs3 ),
       .io_ctrl_mem_ctrl_wfd( ctrl_io_dpath_mem_ctrl_wfd ),
       .io_ctrl_mem_ctrl_div( ctrl_io_dpath_mem_ctrl_div ),
       .io_ctrl_mem_ctrl_wxd( ctrl_io_dpath_mem_ctrl_wxd ),
       .io_ctrl_mem_ctrl_csr( ctrl_io_dpath_mem_ctrl_csr ),
       .io_ctrl_mem_ctrl_fence_i( ctrl_io_dpath_mem_ctrl_fence_i ),
       .io_ctrl_mem_ctrl_sret( ctrl_io_dpath_mem_ctrl_sret ),
       .io_ctrl_mem_ctrl_scall( ctrl_io_dpath_mem_ctrl_scall ),
       .io_ctrl_mem_ctrl_fence( ctrl_io_dpath_mem_ctrl_fence ),
       .io_ctrl_mem_ctrl_amo( ctrl_io_dpath_mem_ctrl_amo ),
       .io_ctrl_csr( ctrl_io_dpath_csr ),
       .io_ctrl_sret( ctrl_io_dpath_sret ),
       .io_ctrl_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_ctrl_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_ctrl_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_ctrl_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_ctrl_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_ctrl_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_ctrl_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_ctrl_retire( ctrl_io_dpath_retire ),
       .io_ctrl_exception( ctrl_io_dpath_exception ),
       .io_ctrl_cause( ctrl_io_dpath_cause ),
       .io_ctrl_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_ctrl_inst( dpath_io_ctrl_inst ),
       .io_ctrl_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_ctrl_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_ctrl_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_ctrl_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_ctrl_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_ctrl_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_ctrl_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_ctrl_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_ctrl_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_ctrl_status_ip( dpath_io_ctrl_status_ip ),
       .io_ctrl_status_im( dpath_io_ctrl_status_im ),
       .io_ctrl_status_zero( dpath_io_ctrl_status_zero ),
       .io_ctrl_status_er( dpath_io_ctrl_status_er ),
       .io_ctrl_status_vm( dpath_io_ctrl_status_vm ),
       .io_ctrl_status_s64( dpath_io_ctrl_status_s64 ),
       .io_ctrl_status_u64( dpath_io_ctrl_status_u64 ),
       .io_ctrl_status_ef( dpath_io_ctrl_status_ef ),
       .io_ctrl_status_pei( dpath_io_ctrl_status_pei ),
       .io_ctrl_status_ei( dpath_io_ctrl_status_ei ),
       .io_ctrl_status_ps( dpath_io_ctrl_status_ps ),
       .io_ctrl_status_s( dpath_io_ctrl_status_s ),
       .io_ctrl_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_ctrl_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_ctrl_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       //.io_dmem_req_valid(  )
       //.io_dmem_req_bits_kill(  )
       //.io_dmem_req_bits_typ(  )
       //.io_dmem_req_bits_phys(  )
       .io_dmem_req_bits_addr( dpath_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( dpath_io_dmem_req_bits_tag ),
       //.io_dmem_req_bits_cmd(  )
       .io_dmem_req_bits_data( dpath_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_ptw_ptbr( dpath_io_ptw_ptbr ),
       .io_ptw_invalidate( dpath_io_ptw_invalidate ),
       .io_ptw_sret( dpath_io_ptw_sret ),
       .io_ptw_status_ip( dpath_io_ptw_status_ip ),
       .io_ptw_status_im( dpath_io_ptw_status_im ),
       .io_ptw_status_zero( dpath_io_ptw_status_zero ),
       .io_ptw_status_er( dpath_io_ptw_status_er ),
       .io_ptw_status_vm( dpath_io_ptw_status_vm ),
       .io_ptw_status_s64( dpath_io_ptw_status_s64 ),
       .io_ptw_status_u64( dpath_io_ptw_status_u64 ),
       .io_ptw_status_ef( dpath_io_ptw_status_ef ),
       .io_ptw_status_pei( dpath_io_ptw_status_pei ),
       .io_ptw_status_ei( dpath_io_ptw_status_ei ),
       .io_ptw_status_ps( dpath_io_ptw_status_ps ),
       .io_ptw_status_s( dpath_io_ptw_status_s ),
       //.io_imem_req_valid(  )
       .io_imem_req_bits_pc( dpath_io_imem_req_bits_pc ),
       //.io_imem_resp_ready(  )
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data_0( io_imem_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( io_imem_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( io_imem_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( io_imem_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( io_imem_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       //.io_imem_btb_update_valid(  )
       //.io_imem_btb_update_bits_prediction_valid(  )
       //.io_imem_btb_update_bits_prediction_bits_taken(  )
       //.io_imem_btb_update_bits_prediction_bits_mask(  )
       //.io_imem_btb_update_bits_prediction_bits_bridx(  )
       //.io_imem_btb_update_bits_prediction_bits_target(  )
       //.io_imem_btb_update_bits_prediction_bits_entry(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_history(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_value(  )
       .io_imem_btb_update_bits_pc( dpath_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( dpath_io_imem_btb_update_bits_target ),
       //.io_imem_btb_update_bits_taken(  )
       //.io_imem_btb_update_bits_isJump(  )
       //.io_imem_btb_update_bits_isReturn(  )
       .io_imem_btb_update_bits_br_pc( dpath_io_imem_btb_update_bits_br_pc ),
       //.io_imem_bht_update_valid(  )
       //.io_imem_bht_update_bits_prediction_valid(  )
       //.io_imem_bht_update_bits_prediction_bits_taken(  )
       //.io_imem_bht_update_bits_prediction_bits_mask(  )
       //.io_imem_bht_update_bits_prediction_bits_bridx(  )
       //.io_imem_bht_update_bits_prediction_bits_target(  )
       //.io_imem_bht_update_bits_prediction_bits_entry(  )
       //.io_imem_bht_update_bits_prediction_bits_bht_history(  )
       //.io_imem_bht_update_bits_prediction_bits_bht_value(  )
       .io_imem_bht_update_bits_pc( dpath_io_imem_bht_update_bits_pc ),
       //.io_imem_bht_update_bits_taken(  )
       //.io_imem_bht_update_bits_mispredict(  )
       //.io_imem_ras_update_valid(  )
       //.io_imem_ras_update_bits_isCall(  )
       //.io_imem_ras_update_bits_isReturn(  )
       .io_imem_ras_update_bits_returnAddr( dpath_io_imem_ras_update_bits_returnAddr ),
       //.io_imem_ras_update_bits_prediction_valid(  )
       //.io_imem_ras_update_bits_prediction_bits_taken(  )
       //.io_imem_ras_update_bits_prediction_bits_mask(  )
       //.io_imem_ras_update_bits_prediction_bits_bridx(  )
       //.io_imem_ras_update_bits_prediction_bits_target(  )
       //.io_imem_ras_update_bits_prediction_bits_entry(  )
       //.io_imem_ras_update_bits_prediction_bits_bht_history(  )
       //.io_imem_ras_update_bits_prediction_bits_bht_value(  )
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       //.io_imem_invalidate(  )
       .io_fpu_inst( dpath_io_fpu_inst ),
       .io_fpu_fromint_data( dpath_io_fpu_fromint_data ),
       .io_fpu_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_fpu_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_fpu_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_fpu_store_data( FPU_io_dpath_store_data ),
       .io_fpu_toint_data( FPU_io_dpath_toint_data ),
       .io_fpu_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_fpu_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_fpu_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_fpu_dmem_resp_data( dpath_io_fpu_dmem_resp_data ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       .io_rocc_cmd_bits_inst_funct( dpath_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( dpath_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( dpath_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( dpath_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( dpath_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( dpath_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( dpath_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( dpath_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( dpath_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( dpath_io_rocc_cmd_bits_rs2 ),
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_uncached( io_rocc_imem_acquire_bits_payload_uncached ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_subblock( io_rocc_imem_acquire_bits_payload_subblock ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_manager_xact_id( io_rocc_imem_finish_bits_payload_manager_xact_id ),
       //.io_rocc_dmem_acquire_ready(  )
       .io_rocc_dmem_acquire_valid( io_rocc_dmem_acquire_valid ),
       .io_rocc_dmem_acquire_bits_header_src( io_rocc_dmem_acquire_bits_header_src ),
       .io_rocc_dmem_acquire_bits_header_dst( io_rocc_dmem_acquire_bits_header_dst ),
       .io_rocc_dmem_acquire_bits_payload_addr( io_rocc_dmem_acquire_bits_payload_addr ),
       .io_rocc_dmem_acquire_bits_payload_client_xact_id( io_rocc_dmem_acquire_bits_payload_client_xact_id ),
       .io_rocc_dmem_acquire_bits_payload_data( io_rocc_dmem_acquire_bits_payload_data ),
       .io_rocc_dmem_acquire_bits_payload_uncached( io_rocc_dmem_acquire_bits_payload_uncached ),
       .io_rocc_dmem_acquire_bits_payload_a_type( io_rocc_dmem_acquire_bits_payload_a_type ),
       .io_rocc_dmem_acquire_bits_payload_subblock( io_rocc_dmem_acquire_bits_payload_subblock ),
       .io_rocc_dmem_grant_ready( io_rocc_dmem_grant_ready ),
       //.io_rocc_dmem_grant_valid(  )
       //.io_rocc_dmem_grant_bits_header_src(  )
       //.io_rocc_dmem_grant_bits_header_dst(  )
       //.io_rocc_dmem_grant_bits_payload_data(  )
       //.io_rocc_dmem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_uncached(  )
       //.io_rocc_dmem_grant_bits_payload_g_type(  )
       //.io_rocc_dmem_finish_ready(  )
       .io_rocc_dmem_finish_valid( io_rocc_dmem_finish_valid ),
       .io_rocc_dmem_finish_bits_header_src( io_rocc_dmem_finish_bits_header_src ),
       .io_rocc_dmem_finish_bits_header_dst( io_rocc_dmem_finish_bits_header_dst ),
       .io_rocc_dmem_finish_bits_payload_manager_xact_id( io_rocc_dmem_finish_bits_payload_manager_xact_id ),
       .io_rocc_dmem_probe_ready( io_rocc_dmem_probe_ready ),
       //.io_rocc_dmem_probe_valid(  )
       //.io_rocc_dmem_probe_bits_header_src(  )
       //.io_rocc_dmem_probe_bits_header_dst(  )
       //.io_rocc_dmem_probe_bits_payload_addr(  )
       //.io_rocc_dmem_probe_bits_payload_p_type(  )
       //.io_rocc_dmem_release_ready(  )
       .io_rocc_dmem_release_valid( io_rocc_dmem_release_valid ),
       .io_rocc_dmem_release_bits_header_src( io_rocc_dmem_release_bits_header_src ),
       .io_rocc_dmem_release_bits_header_dst( io_rocc_dmem_release_bits_header_dst ),
       .io_rocc_dmem_release_bits_payload_addr( io_rocc_dmem_release_bits_payload_addr ),
       .io_rocc_dmem_release_bits_payload_client_xact_id( io_rocc_dmem_release_bits_payload_client_xact_id ),
       .io_rocc_dmem_release_bits_payload_data( io_rocc_dmem_release_bits_payload_data ),
       .io_rocc_dmem_release_bits_payload_r_type( io_rocc_dmem_release_bits_payload_r_type ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  FPU FPU(.clk(clk), .reset(reset),
       .io_ctrl_valid( ctrl_io_fpu_valid ),
       .io_ctrl_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_ctrl_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_ctrl_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_ctrl_killx( ctrl_io_fpu_killx ),
       .io_ctrl_killm( ctrl_io_fpu_killm ),
       .io_ctrl_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_ctrl_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_ctrl_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_ctrl_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_ctrl_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_ctrl_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_ctrl_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_ctrl_dec_single( FPU_io_ctrl_dec_single ),
       .io_ctrl_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_ctrl_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_ctrl_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_ctrl_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_ctrl_dec_round( FPU_io_ctrl_dec_round ),
       .io_ctrl_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_ctrl_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_ctrl_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_dpath_inst( dpath_io_fpu_inst ),
       .io_dpath_fromint_data( dpath_io_fpu_fromint_data ),
       .io_dpath_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_dpath_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_dpath_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_dpath_store_data( FPU_io_dpath_store_data ),
       .io_dpath_toint_data( FPU_io_dpath_toint_data ),
       .io_dpath_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_dpath_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_dpath_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_dpath_dmem_resp_data( dpath_io_fpu_dmem_resp_data )
  );
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input  io_requestor_1_req_bits_kill,
    input [3:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_phys,
    input [43:0] io_requestor_1_req_bits_addr,
    input [7:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    input [63:0] io_requestor_1_req_bits_data,
    output io_requestor_1_resp_valid,
    output[63:0] io_requestor_1_resp_bits_data,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output[3:0] io_requestor_1_resp_bits_typ,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[7:0] io_requestor_1_resp_bits_tag,
    output[3:0] io_requestor_1_resp_bits_cmd,
    output[43:0] io_requestor_1_resp_bits_addr,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[7:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    //input  io_requestor_1_ptw_req_ready
    //output io_requestor_1_ptw_req_valid
    //output[29:0] io_requestor_1_ptw_req_bits
    //input  io_requestor_1_ptw_resp_valid
    //input  io_requestor_1_ptw_resp_bits_error
    //input [18:0] io_requestor_1_ptw_resp_bits_ppn
    //input [5:0] io_requestor_1_ptw_resp_bits_perm
    //input [7:0] io_requestor_1_ptw_status_ip
    //input [7:0] io_requestor_1_ptw_status_im
    //input [6:0] io_requestor_1_ptw_status_zero
    //input  io_requestor_1_ptw_status_er
    //input  io_requestor_1_ptw_status_vm
    //input  io_requestor_1_ptw_status_s64
    //input  io_requestor_1_ptw_status_u64
    //input  io_requestor_1_ptw_status_ef
    //input  io_requestor_1_ptw_status_pei
    //input  io_requestor_1_ptw_status_ei
    //input  io_requestor_1_ptw_status_ps
    //input  io_requestor_1_ptw_status_s
    //input  io_requestor_1_ptw_invalidate
    //input  io_requestor_1_ptw_sret
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input  io_requestor_0_req_bits_kill,
    input [3:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_phys,
    input [43:0] io_requestor_0_req_bits_addr,
    input [7:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    input [63:0] io_requestor_0_req_bits_data,
    output io_requestor_0_resp_valid,
    output[63:0] io_requestor_0_resp_bits_data,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output[3:0] io_requestor_0_resp_bits_typ,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[7:0] io_requestor_0_resp_bits_tag,
    output[3:0] io_requestor_0_resp_bits_cmd,
    output[43:0] io_requestor_0_resp_bits_addr,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[7:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_ptw_req_ready
    //output io_requestor_0_ptw_req_valid
    //output[29:0] io_requestor_0_ptw_req_bits
    //input  io_requestor_0_ptw_resp_valid
    //input  io_requestor_0_ptw_resp_bits_error
    //input [18:0] io_requestor_0_ptw_resp_bits_ppn
    //input [5:0] io_requestor_0_ptw_resp_bits_perm
    //input [7:0] io_requestor_0_ptw_status_ip
    //input [7:0] io_requestor_0_ptw_status_im
    //input [6:0] io_requestor_0_ptw_status_zero
    //input  io_requestor_0_ptw_status_er
    //input  io_requestor_0_ptw_status_vm
    //input  io_requestor_0_ptw_status_s64
    //input  io_requestor_0_ptw_status_u64
    //input  io_requestor_0_ptw_status_ef
    //input  io_requestor_0_ptw_status_pei
    //input  io_requestor_0_ptw_status_ei
    //input  io_requestor_0_ptw_status_ps
    //input  io_requestor_0_ptw_status_s
    //input  io_requestor_0_ptw_invalidate
    //input  io_requestor_0_ptw_sret
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[3:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    output[7:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [3:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered
);

  wire[63:0] T0;
  reg  r_valid_0;
  wire[4:0] T1;
  wire[7:0] T32;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[8:0] T4;
  wire[43:0] T5;
  wire T6;
  wire[3:0] T7;
  wire T8;
  wire T9;
  wire[7:0] T33;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[7:0] T34;
  wire[6:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[7:0] T35;
  wire[6:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[7:0] T36;
  wire[6:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
// synthesis translate_on
`endif

//  assign io_mem_ptw_sret = {1{$random}};
//  assign io_mem_ptw_invalidate = {1{$random}};
//  assign io_mem_ptw_status_s = {1{$random}};
//  assign io_mem_ptw_status_ps = {1{$random}};
//  assign io_mem_ptw_status_ei = {1{$random}};
//  assign io_mem_ptw_status_pei = {1{$random}};
//  assign io_mem_ptw_status_ef = {1{$random}};
//  assign io_mem_ptw_status_u64 = {1{$random}};
//  assign io_mem_ptw_status_s64 = {1{$random}};
//  assign io_mem_ptw_status_vm = {1{$random}};
//  assign io_mem_ptw_status_er = {1{$random}};
//  assign io_mem_ptw_status_zero = {1{$random}};
//  assign io_mem_ptw_status_im = {1{$random}};
//  assign io_mem_ptw_status_ip = {1{$random}};
//  assign io_mem_ptw_resp_bits_perm = {1{$random}};
//  assign io_mem_ptw_resp_bits_ppn = {1{$random}};
//  assign io_mem_ptw_resp_bits_error = {1{$random}};
//  assign io_mem_ptw_resp_valid = {1{$random}};
//  assign io_mem_ptw_req_ready = {1{$random}};
  assign io_mem_req_bits_data = T0;
  assign T0 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_cmd = T1;
  assign T1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T32;
  assign T32 = T2[3'h7:1'h0];
  assign T2 = io_requestor_0_req_valid ? T4 : T3;
  assign T3 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T4 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_addr = T5;
  assign T5 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_bits_phys = T6;
  assign T6 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_typ = T7;
  assign T7 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_kill = T8;
  assign T8 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_valid = T9;
  assign T9 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
//  assign io_requestor_0_ptw_req_bits = {1{$random}};
//  assign io_requestor_0_ptw_req_valid = {1{$random}};
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T33;
  assign T33 = {1'h0, T10};
  assign T10 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T11;
  assign T11 = io_mem_replay_next_valid & T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T34;
  assign T34 = {1'h0, T14};
  assign T14 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_replay = T15;
  assign T15 = io_mem_resp_bits_replay & T16;
  assign T16 = T17 == 1'h0;
  assign T17 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T18;
  assign T18 = io_mem_resp_bits_nack & T16;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_valid = T19;
  assign T19 = io_mem_resp_valid & T16;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
//  assign io_requestor_1_ptw_req_bits = {1{$random}};
//  assign io_requestor_1_ptw_req_valid = {1{$random}};
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T35;
  assign T35 = {1'h0, T20};
  assign T20 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T21;
  assign T21 = io_mem_replay_next_valid & T22;
  assign T22 = T23 == 1'h1;
  assign T23 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T36;
  assign T36 = {1'h0, T24};
  assign T24 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_replay = T25;
  assign T25 = io_mem_resp_bits_replay & T26;
  assign T26 = T27 == 1'h1;
  assign T27 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T28;
  assign T28 = io_mem_resp_bits_nack & T26;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_valid = T29;
  assign T29 = io_mem_resp_valid & T26;
  assign io_requestor_1_req_ready = T30;
  assign T30 = io_requestor_0_req_ready & T31;
  assign T31 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [135:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [128:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [135:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [128:0] io_in_0_bits_payload_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[135:0] io_out_bits_payload_data,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_a_type,
    output[128:0] io_out_bits_payload_subblock,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T55;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T56;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg  locked;
  wire T57;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] T21;
  reg [1:0] R22;
  wire[1:0] T58;
  wire[1:0] T23;
  wire[128:0] T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire[135:0] T28;
  wire[1:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R22 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T55 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T56 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T16 & T12;
  assign T12 = io_out_bits_payload_uncached ? T13 : 1'h0;
  assign T13 = T15 | T14;
  assign T14 = 2'h2 == io_out_bits_payload_a_type;
  assign T15 = 2'h1 == io_out_bits_payload_a_type;
  assign T16 = io_out_ready & io_out_valid;
  assign T57 = reset ? 1'h0 : T17;
  assign T17 = T19 ? 1'h0 : T18;
  assign T18 = T9 ? 1'h1 : locked;
  assign T19 = T16 & T20;
  assign T20 = T21 == 2'h0;
  assign T21 = R22 + 2'h1;
  assign T58 = reset ? 2'h0 : T23;
  assign T23 = T11 ? T21 : R22;
  assign io_out_bits_payload_subblock = T24;
  assign T24 = T25 ? io_in_1_bits_payload_subblock : io_in_0_bits_payload_subblock;
  assign T25 = chosen;
  assign io_out_bits_payload_a_type = T26;
  assign T26 = T25 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign io_out_bits_payload_uncached = T27;
  assign T27 = T25 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign io_out_bits_payload_data = T28;
  assign T28 = T25 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign io_out_bits_payload_client_xact_id = T29;
  assign T29 = T25 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr = T30;
  assign T30 = T25 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign io_out_bits_header_dst = T31;
  assign T31 = T25 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T32;
  assign T32 = T25 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T33;
  assign T33 = T25 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T34;
  assign T34 = T35 & io_out_ready;
  assign T35 = locked ? T44 : T36;
  assign T36 = T43 | T37;
  assign T37 = T38 ^ 1'h1;
  assign T38 = T41 | T39;
  assign T39 = io_in_1_valid & T40;
  assign T40 = last_grant < 1'h1;
  assign T41 = io_in_0_valid & T42;
  assign T42 = last_grant < 1'h0;
  assign T43 = last_grant < 1'h0;
  assign T44 = lockIdx == 1'h0;
  assign io_in_1_ready = T45;
  assign T45 = T46 & io_out_ready;
  assign T46 = locked ? T54 : T47;
  assign T47 = T51 | T48;
  assign T48 = T49 ^ 1'h1;
  assign T49 = T50 | io_in_0_valid;
  assign T50 = T41 | T39;
  assign T51 = T53 & T52;
  assign T52 = last_grant < 1'h1;
  assign T53 = T41 ^ 1'h1;
  assign T54 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T19) begin
      locked <= 1'h0;
    end else if(T9) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R22 <= 2'h0;
    end else if(T11) begin
      R22 <= T21;
    end
  end
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [135:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [135:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[135:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T56;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T57;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg  locked;
  wire T58;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  reg [1:0] R25;
  wire[1:0] T59;
  wire[1:0] T26;
  wire[2:0] T27;
  wire T28;
  wire[135:0] T29;
  wire[1:0] T30;
  wire[25:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R25 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T56 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T57 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T19 & T12;
  assign T12 = T14 | T13;
  assign T13 = 3'h3 == io_out_bits_payload_r_type;
  assign T14 = T16 | T15;
  assign T15 = 3'h2 == io_out_bits_payload_r_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h1 == io_out_bits_payload_r_type;
  assign T18 = 3'h0 == io_out_bits_payload_r_type;
  assign T19 = io_out_ready & io_out_valid;
  assign T58 = reset ? 1'h0 : T20;
  assign T20 = T22 ? 1'h0 : T21;
  assign T21 = T9 ? 1'h1 : locked;
  assign T22 = T19 & T23;
  assign T23 = T24 == 2'h0;
  assign T24 = R25 + 2'h1;
  assign T59 = reset ? 2'h0 : T26;
  assign T26 = T11 ? T24 : R25;
  assign io_out_bits_payload_r_type = T27;
  assign T27 = T28 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T28 = chosen;
  assign io_out_bits_payload_data = T29;
  assign T29 = T28 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign io_out_bits_payload_client_xact_id = T30;
  assign T30 = T28 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr = T31;
  assign T31 = T28 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign io_out_bits_header_dst = T32;
  assign T32 = T28 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T33;
  assign T33 = T28 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T34;
  assign T34 = T28 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T35;
  assign T35 = T36 & io_out_ready;
  assign T36 = locked ? T45 : T37;
  assign T37 = T44 | T38;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T42 | T40;
  assign T40 = io_in_1_valid & T41;
  assign T41 = last_grant < 1'h1;
  assign T42 = io_in_0_valid & T43;
  assign T43 = last_grant < 1'h0;
  assign T44 = last_grant < 1'h0;
  assign T45 = lockIdx == 1'h0;
  assign io_in_1_ready = T46;
  assign T46 = T47 & io_out_ready;
  assign T47 = locked ? T55 : T48;
  assign T48 = T52 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_0_valid;
  assign T51 = T42 | T40;
  assign T52 = T54 & T53;
  assign T53 = last_grant < 1'h1;
  assign T54 = T42 ^ 1'h1;
  assign T55 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T22) begin
      locked <= 1'h0;
    end else if(T9) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R25 <= 2'h0;
    end else if(T11) begin
      R25 <= T24;
    end
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[3:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_manager_xact_id = T5;
  assign T5 = T6 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T6 = chosen;
  assign io_out_bits_header_dst = T7;
  assign T7 = T6 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T8;
  assign T8 = T6 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module TileLinkIOArbiterThatAppendsArbiterId(input clk, input reset,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [1:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [135:0] io_in_1_acquire_bits_payload_data,
    input  io_in_1_acquire_bits_payload_uncached,
    input [1:0] io_in_1_acquire_bits_payload_a_type,
    input [128:0] io_in_1_acquire_bits_payload_subblock,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[135:0] io_in_1_grant_bits_payload_data,
    output[1:0] io_in_1_grant_bits_payload_client_xact_id,
    output[3:0] io_in_1_grant_bits_payload_manager_xact_id,
    output io_in_1_grant_bits_payload_uncached,
    output[1:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [3:0] io_in_1_finish_bits_payload_manager_xact_id,
    input  io_in_1_probe_ready,
    output io_in_1_probe_valid,
    output[1:0] io_in_1_probe_bits_header_src,
    output[1:0] io_in_1_probe_bits_header_dst,
    output[25:0] io_in_1_probe_bits_payload_addr,
    output[1:0] io_in_1_probe_bits_payload_p_type,
    output io_in_1_release_ready,
    input  io_in_1_release_valid,
    input [1:0] io_in_1_release_bits_header_src,
    input [1:0] io_in_1_release_bits_header_dst,
    input [25:0] io_in_1_release_bits_payload_addr,
    input [1:0] io_in_1_release_bits_payload_client_xact_id,
    input [135:0] io_in_1_release_bits_payload_data,
    input [2:0] io_in_1_release_bits_payload_r_type,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [1:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [135:0] io_in_0_acquire_bits_payload_data,
    input  io_in_0_acquire_bits_payload_uncached,
    input [1:0] io_in_0_acquire_bits_payload_a_type,
    input [128:0] io_in_0_acquire_bits_payload_subblock,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[135:0] io_in_0_grant_bits_payload_data,
    output[1:0] io_in_0_grant_bits_payload_client_xact_id,
    output[3:0] io_in_0_grant_bits_payload_manager_xact_id,
    output io_in_0_grant_bits_payload_uncached,
    output[1:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [3:0] io_in_0_finish_bits_payload_manager_xact_id,
    input  io_in_0_probe_ready,
    output io_in_0_probe_valid,
    output[1:0] io_in_0_probe_bits_header_src,
    output[1:0] io_in_0_probe_bits_header_dst,
    output[25:0] io_in_0_probe_bits_payload_addr,
    output[1:0] io_in_0_probe_bits_payload_p_type,
    output io_in_0_release_ready,
    input  io_in_0_release_valid,
    input [1:0] io_in_0_release_bits_header_src,
    input [1:0] io_in_0_release_bits_header_dst,
    input [25:0] io_in_0_release_bits_payload_addr,
    input [1:0] io_in_0_release_bits_payload_client_xact_id,
    input [135:0] io_in_0_release_bits_payload_data,
    input [2:0] io_in_0_release_bits_payload_r_type,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[135:0] io_out_acquire_bits_payload_data,
    output io_out_acquire_bits_payload_uncached,
    output[1:0] io_out_acquire_bits_payload_a_type,
    output[128:0] io_out_acquire_bits_payload_subblock,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [135:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [3:0] io_out_grant_bits_payload_manager_xact_id,
    input  io_out_grant_bits_payload_uncached,
    input [1:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[3:0] io_out_finish_bits_payload_manager_xact_id,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [1:0] io_out_probe_bits_header_src,
    input [1:0] io_out_probe_bits_header_dst,
    input [25:0] io_out_probe_bits_payload_addr,
    input [1:0] io_out_probe_bits_payload_p_type,
    input  io_out_release_ready,
    output io_out_release_valid,
    output[1:0] io_out_release_bits_header_src,
    output[1:0] io_out_release_bits_header_dst,
    output[25:0] io_out_release_bits_payload_addr,
    output[1:0] io_out_release_bits_payload_client_xact_id,
    output[135:0] io_out_release_bits_payload_data,
    output[2:0] io_out_release_bits_payload_r_type
);

  wire[1:0] T17;
  wire[2:0] T0;
  wire[1:0] T18;
  wire[2:0] T1;
  wire[1:0] T19;
  wire[2:0] T2;
  wire[1:0] T20;
  wire[2:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire[1:0] T21;
  wire T13;
  wire T14;
  wire[1:0] T22;
  wire T15;
  wire T16;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire LockingRRArbiter_0_io_out_valid;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire LockingRRArbiter_0_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_a_type;
  wire[128:0] LockingRRArbiter_0_io_out_bits_payload_subblock;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire finish_arb_io_in_1_ready;
  wire finish_arb_io_in_0_ready;
  wire finish_arb_io_out_valid;
  wire[1:0] finish_arb_io_out_bits_header_src;
  wire[1:0] finish_arb_io_out_bits_header_dst;
  wire[3:0] finish_arb_io_out_bits_payload_manager_xact_id;


  assign T17 = T0[1'h1:1'h0];
  assign T0 = {io_in_0_release_bits_payload_client_xact_id, 1'h0};
  assign T18 = T1[1'h1:1'h0];
  assign T1 = {io_in_1_release_bits_payload_client_xact_id, 1'h1};
  assign T19 = T2[1'h1:1'h0];
  assign T2 = {io_in_0_acquire_bits_payload_client_xact_id, 1'h0};
  assign T20 = T3[1'h1:1'h0];
  assign T3 = {io_in_1_acquire_bits_payload_client_xact_id, 1'h1};
  assign io_out_release_bits_payload_r_type = LockingRRArbiter_1_io_out_bits_payload_r_type;
  assign io_out_release_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_release_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_release_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_release_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_release_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_release_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_probe_ready = T4;
  assign T4 = io_in_0_probe_ready | io_in_1_probe_ready;
  assign io_out_finish_bits_payload_manager_xact_id = finish_arb_io_out_bits_payload_manager_xact_id;
  assign io_out_finish_bits_header_dst = finish_arb_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = finish_arb_io_out_bits_header_src;
  assign io_out_finish_valid = finish_arb_io_out_valid;
  assign io_out_grant_ready = T5;
  assign T5 = T10 ? io_in_1_grant_ready : T6;
  assign T6 = T7 ? io_in_0_grant_ready : 1'h0;
  assign T7 = T8 == 1'h0;
  assign T8 = T9;
  assign T9 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign T10 = T11 == 1'h1;
  assign T11 = T12;
  assign T12 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_out_acquire_bits_payload_subblock = LockingRRArbiter_0_io_out_bits_payload_subblock;
  assign io_out_acquire_bits_payload_a_type = LockingRRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_uncached = LockingRRArbiter_0_io_out_bits_payload_uncached;
  assign io_out_acquire_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = LockingRRArbiter_0_io_out_valid;
  assign io_in_0_release_ready = LockingRRArbiter_1_io_in_0_ready;
  assign io_in_0_probe_bits_payload_p_type = io_out_probe_bits_payload_p_type;
  assign io_in_0_probe_bits_payload_addr = io_out_probe_bits_payload_addr;
  assign io_in_0_probe_bits_header_dst = io_out_probe_bits_header_dst;
  assign io_in_0_probe_bits_header_src = io_out_probe_bits_header_src;
  assign io_in_0_probe_valid = io_out_probe_valid;
  assign io_in_0_finish_ready = finish_arb_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_0_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = T21;
  assign T21 = {1'h0, T13};
  assign T13 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T14;
  assign T14 = T7 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_0_io_in_0_ready;
  assign io_in_1_release_ready = LockingRRArbiter_1_io_in_1_ready;
  assign io_in_1_probe_bits_payload_p_type = io_out_probe_bits_payload_p_type;
  assign io_in_1_probe_bits_payload_addr = io_out_probe_bits_payload_addr;
  assign io_in_1_probe_bits_header_dst = io_out_probe_bits_header_dst;
  assign io_in_1_probe_bits_header_src = io_out_probe_bits_header_src;
  assign io_in_1_probe_valid = io_out_probe_valid;
  assign io_in_1_finish_ready = finish_arb_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_1_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = T22;
  assign T22 = {1'h0, T15};
  assign T15 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T16;
  assign T16 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_0_io_in_1_ready;
  LockingRRArbiter_0 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T20 ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_acquire_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_acquire_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T19 ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_acquire_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_acquire_bits_payload_subblock ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_0_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_0_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_release_valid ),
       .io_in_1_bits_header_src( io_in_1_release_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_release_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_release_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T18 ),
       .io_in_1_bits_payload_data( io_in_1_release_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_release_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_release_valid ),
       .io_in_0_bits_header_src( io_in_0_release_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_release_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_release_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T17 ),
       .io_in_0_bits_payload_data( io_in_0_release_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_release_bits_payload_r_type ),
       .io_out_ready( io_out_release_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  RRArbiter_1 finish_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( finish_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_finish_bits_payload_manager_xact_id ),
       .io_in_0_ready( finish_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_finish_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( finish_arb_io_out_valid ),
       .io_out_bits_header_src( finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( finish_arb_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module TileLinkIOWrapper(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [1:0] io_in_acquire_bits_header_src,
    input [1:0] io_in_acquire_bits_header_dst,
    input [25:0] io_in_acquire_bits_payload_addr,
    input [1:0] io_in_acquire_bits_payload_client_xact_id,
    input [135:0] io_in_acquire_bits_payload_data,
    input  io_in_acquire_bits_payload_uncached,
    input [1:0] io_in_acquire_bits_payload_a_type,
    input [128:0] io_in_acquire_bits_payload_subblock,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_header_src,
    output[1:0] io_in_grant_bits_header_dst,
    output[135:0] io_in_grant_bits_payload_data,
    output[1:0] io_in_grant_bits_payload_client_xact_id,
    output[3:0] io_in_grant_bits_payload_manager_xact_id,
    output io_in_grant_bits_payload_uncached,
    output[1:0] io_in_grant_bits_payload_g_type,
    output io_in_finish_ready,
    input  io_in_finish_valid,
    input [1:0] io_in_finish_bits_header_src,
    input [1:0] io_in_finish_bits_header_dst,
    input [3:0] io_in_finish_bits_payload_manager_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[135:0] io_out_acquire_bits_payload_data,
    output io_out_acquire_bits_payload_uncached,
    output[1:0] io_out_acquire_bits_payload_a_type,
    output[128:0] io_out_acquire_bits_payload_subblock,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [135:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [3:0] io_out_grant_bits_payload_manager_xact_id,
    input  io_out_grant_bits_payload_uncached,
    input [1:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[3:0] io_out_finish_bits_payload_manager_xact_id,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [1:0] io_out_probe_bits_header_src,
    input [1:0] io_out_probe_bits_header_dst,
    input [25:0] io_out_probe_bits_payload_addr,
    input [1:0] io_out_probe_bits_payload_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_header_src
    //output[1:0] io_out_release_bits_header_dst
    //output[25:0] io_out_release_bits_payload_addr
    //output[1:0] io_out_release_bits_payload_client_xact_id
    //output[135:0] io_out_release_bits_payload_data
    //output[2:0] io_out_release_bits_payload_r_type
);



//  assign io_out_release_bits_payload_r_type = {1{$random}};
//  assign io_out_release_bits_payload_data = {5{$random}};
//  assign io_out_release_bits_payload_client_xact_id = {1{$random}};
//  assign io_out_release_bits_payload_addr = {1{$random}};
//  assign io_out_release_bits_header_dst = {1{$random}};
//  assign io_out_release_bits_header_src = {1{$random}};
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h0;
  assign io_out_finish_bits_payload_manager_xact_id = io_in_finish_bits_payload_manager_xact_id;
  assign io_out_finish_bits_header_dst = io_in_finish_bits_header_dst;
  assign io_out_finish_bits_header_src = io_in_finish_bits_header_src;
  assign io_out_finish_valid = io_in_finish_valid;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_payload_subblock = io_in_acquire_bits_payload_subblock;
  assign io_out_acquire_bits_payload_a_type = io_in_acquire_bits_payload_a_type;
  assign io_out_acquire_bits_payload_uncached = io_in_acquire_bits_payload_uncached;
  assign io_out_acquire_bits_payload_data = io_in_acquire_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = io_in_acquire_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = io_in_acquire_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = io_in_acquire_bits_header_dst;
  assign io_out_acquire_bits_header_src = io_in_acquire_bits_header_src;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_finish_ready = io_out_finish_ready;
  assign io_in_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module RocketTile(input clk, input reset,
    input  io_tilelink_acquire_ready,
    output io_tilelink_acquire_valid,
    output[1:0] io_tilelink_acquire_bits_header_src,
    output[1:0] io_tilelink_acquire_bits_header_dst,
    output[25:0] io_tilelink_acquire_bits_payload_addr,
    output[1:0] io_tilelink_acquire_bits_payload_client_xact_id,
    output[135:0] io_tilelink_acquire_bits_payload_data,
    output io_tilelink_acquire_bits_payload_uncached,
    output[1:0] io_tilelink_acquire_bits_payload_a_type,
    output[128:0] io_tilelink_acquire_bits_payload_subblock,
    output io_tilelink_grant_ready,
    input  io_tilelink_grant_valid,
    input [1:0] io_tilelink_grant_bits_header_src,
    input [1:0] io_tilelink_grant_bits_header_dst,
    input [135:0] io_tilelink_grant_bits_payload_data,
    input [1:0] io_tilelink_grant_bits_payload_client_xact_id,
    input [3:0] io_tilelink_grant_bits_payload_manager_xact_id,
    input  io_tilelink_grant_bits_payload_uncached,
    input [1:0] io_tilelink_grant_bits_payload_g_type,
    input  io_tilelink_finish_ready,
    output io_tilelink_finish_valid,
    output[1:0] io_tilelink_finish_bits_header_src,
    output[1:0] io_tilelink_finish_bits_header_dst,
    output[3:0] io_tilelink_finish_bits_payload_manager_xact_id,
    output io_tilelink_probe_ready,
    input  io_tilelink_probe_valid,
    input [1:0] io_tilelink_probe_bits_header_src,
    input [1:0] io_tilelink_probe_bits_header_dst,
    input [25:0] io_tilelink_probe_bits_payload_addr,
    input [1:0] io_tilelink_probe_bits_payload_p_type,
    input  io_tilelink_release_ready,
    output io_tilelink_release_valid,
    output[1:0] io_tilelink_release_bits_header_src,
    output[1:0] io_tilelink_release_bits_header_dst,
    output[25:0] io_tilelink_release_bits_payload_addr,
    output[1:0] io_tilelink_release_bits_payload_client_xact_id,
    output[135:0] io_tilelink_release_bits_payload_data,
    output[2:0] io_tilelink_release_bits_payload_r_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr
);

  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire[3:0] dcArb_io_requestor_1_resp_bits_typ;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_subword;
  wire[7:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[7:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire[3:0] dcArb_io_requestor_0_resp_bits_typ;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_subword;
  wire[7:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[7:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire dcArb_io_mem_req_bits_kill;
  wire[3:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_phys;
  wire[43:0] dcArb_io_mem_req_bits_addr;
  wire[7:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire TileLinkIOWrapper_io_in_acquire_ready;
  wire TileLinkIOWrapper_io_in_grant_valid;
  wire[1:0] TileLinkIOWrapper_io_in_grant_bits_header_src;
  wire[1:0] TileLinkIOWrapper_io_in_grant_bits_header_dst;
  wire[135:0] TileLinkIOWrapper_io_in_grant_bits_payload_data;
  wire[1:0] TileLinkIOWrapper_io_in_grant_bits_payload_client_xact_id;
  wire[3:0] TileLinkIOWrapper_io_in_grant_bits_payload_manager_xact_id;
  wire TileLinkIOWrapper_io_in_grant_bits_payload_uncached;
  wire[1:0] TileLinkIOWrapper_io_in_grant_bits_payload_g_type;
  wire TileLinkIOWrapper_io_in_finish_ready;
  wire TileLinkIOWrapper_io_out_acquire_valid;
  wire[1:0] TileLinkIOWrapper_io_out_acquire_bits_header_src;
  wire[1:0] TileLinkIOWrapper_io_out_acquire_bits_header_dst;
  wire[25:0] TileLinkIOWrapper_io_out_acquire_bits_payload_addr;
  wire[1:0] TileLinkIOWrapper_io_out_acquire_bits_payload_client_xact_id;
  wire[135:0] TileLinkIOWrapper_io_out_acquire_bits_payload_data;
  wire TileLinkIOWrapper_io_out_acquire_bits_payload_uncached;
  wire[1:0] TileLinkIOWrapper_io_out_acquire_bits_payload_a_type;
  wire[128:0] TileLinkIOWrapper_io_out_acquire_bits_payload_subblock;
  wire TileLinkIOWrapper_io_out_grant_ready;
  wire TileLinkIOWrapper_io_out_finish_valid;
  wire[1:0] TileLinkIOWrapper_io_out_finish_bits_header_src;
  wire[1:0] TileLinkIOWrapper_io_out_finish_bits_header_dst;
  wire[3:0] TileLinkIOWrapper_io_out_finish_bits_payload_manager_xact_id;
  wire TileLinkIOWrapper_io_out_probe_ready;
  wire TileLinkIOWrapper_io_out_release_valid;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[18:0] ptw_io_requestor_1_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_1_resp_bits_perm;
  wire[7:0] ptw_io_requestor_1_status_ip;
  wire[7:0] ptw_io_requestor_1_status_im;
  wire[6:0] ptw_io_requestor_1_status_zero;
  wire ptw_io_requestor_1_status_er;
  wire ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_s64;
  wire ptw_io_requestor_1_status_u64;
  wire ptw_io_requestor_1_status_ef;
  wire ptw_io_requestor_1_status_pei;
  wire ptw_io_requestor_1_status_ei;
  wire ptw_io_requestor_1_status_ps;
  wire ptw_io_requestor_1_status_s;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_1_sret;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[18:0] ptw_io_requestor_0_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_0_resp_bits_perm;
  wire[7:0] ptw_io_requestor_0_status_ip;
  wire[7:0] ptw_io_requestor_0_status_im;
  wire[6:0] ptw_io_requestor_0_status_zero;
  wire ptw_io_requestor_0_status_er;
  wire ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_s64;
  wire ptw_io_requestor_0_status_u64;
  wire ptw_io_requestor_0_status_ef;
  wire ptw_io_requestor_0_status_pei;
  wire ptw_io_requestor_0_status_ei;
  wire ptw_io_requestor_0_status_ps;
  wire ptw_io_requestor_0_status_s;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_requestor_0_sret;
  wire ptw_io_mem_req_valid;
  wire ptw_io_mem_req_bits_kill;
  wire[3:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_phys;
  wire[43:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire memArb_io_in_1_acquire_ready;
  wire memArb_io_in_1_grant_valid;
  wire[1:0] memArb_io_in_1_grant_bits_header_src;
  wire[1:0] memArb_io_in_1_grant_bits_header_dst;
  wire[135:0] memArb_io_in_1_grant_bits_payload_data;
  wire[1:0] memArb_io_in_1_grant_bits_payload_client_xact_id;
  wire[3:0] memArb_io_in_1_grant_bits_payload_manager_xact_id;
  wire memArb_io_in_1_grant_bits_payload_uncached;
  wire[1:0] memArb_io_in_1_grant_bits_payload_g_type;
  wire memArb_io_in_1_finish_ready;
  wire memArb_io_in_1_probe_valid;
  wire[1:0] memArb_io_in_1_probe_bits_header_src;
  wire[1:0] memArb_io_in_1_probe_bits_header_dst;
  wire[25:0] memArb_io_in_1_probe_bits_payload_addr;
  wire[1:0] memArb_io_in_1_probe_bits_payload_p_type;
  wire memArb_io_in_1_release_ready;
  wire memArb_io_in_0_acquire_ready;
  wire memArb_io_in_0_grant_valid;
  wire[1:0] memArb_io_in_0_grant_bits_header_src;
  wire[1:0] memArb_io_in_0_grant_bits_header_dst;
  wire[135:0] memArb_io_in_0_grant_bits_payload_data;
  wire[1:0] memArb_io_in_0_grant_bits_payload_client_xact_id;
  wire[3:0] memArb_io_in_0_grant_bits_payload_manager_xact_id;
  wire memArb_io_in_0_grant_bits_payload_uncached;
  wire[1:0] memArb_io_in_0_grant_bits_payload_g_type;
  wire memArb_io_in_0_finish_ready;
  wire memArb_io_in_0_probe_valid;
  wire[1:0] memArb_io_in_0_probe_bits_header_src;
  wire[1:0] memArb_io_in_0_probe_bits_header_dst;
  wire[25:0] memArb_io_in_0_probe_bits_payload_addr;
  wire[1:0] memArb_io_in_0_probe_bits_payload_p_type;
  wire memArb_io_in_0_release_ready;
  wire memArb_io_out_acquire_valid;
  wire[1:0] memArb_io_out_acquire_bits_header_src;
  wire[1:0] memArb_io_out_acquire_bits_header_dst;
  wire[25:0] memArb_io_out_acquire_bits_payload_addr;
  wire[1:0] memArb_io_out_acquire_bits_payload_client_xact_id;
  wire[135:0] memArb_io_out_acquire_bits_payload_data;
  wire memArb_io_out_acquire_bits_payload_uncached;
  wire[1:0] memArb_io_out_acquire_bits_payload_a_type;
  wire[128:0] memArb_io_out_acquire_bits_payload_subblock;
  wire memArb_io_out_grant_ready;
  wire memArb_io_out_finish_valid;
  wire[1:0] memArb_io_out_finish_bits_header_src;
  wire[1:0] memArb_io_out_finish_bits_header_dst;
  wire[3:0] memArb_io_out_finish_bits_payload_manager_xact_id;
  wire memArb_io_out_probe_ready;
  wire memArb_io_out_release_valid;
  wire[1:0] memArb_io_out_release_bits_header_src;
  wire[1:0] memArb_io_out_release_bits_header_dst;
  wire[25:0] memArb_io_out_release_bits_payload_addr;
  wire[1:0] memArb_io_out_release_bits_payload_client_xact_id;
  wire[135:0] memArb_io_out_release_bits_payload_data;
  wire[2:0] memArb_io_out_release_bits_payload_r_type;
  wire icache_io_cpu_resp_valid;
  wire[43:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data_0;
  wire icache_io_cpu_resp_bits_mask;
  wire icache_io_cpu_resp_bits_xcpt_ma;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_bits_mask;
  wire icache_io_cpu_btb_resp_bits_bridx;
  wire[42:0] icache_io_cpu_btb_resp_bits_target;
  wire[5:0] icache_io_cpu_btb_resp_bits_entry;
  wire[6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire icache_io_cpu_ptw_req_valid;
  wire[29:0] icache_io_cpu_ptw_req_bits;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[135:0] icache_io_mem_acquire_bits_payload_data;
  wire icache_io_mem_acquire_bits_payload_uncached;
  wire[1:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[128:0] icache_io_mem_acquire_bits_payload_subblock;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[3:0] icache_io_mem_finish_bits_payload_manager_xact_id;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire[3:0] dcache_io_cpu_resp_bits_typ;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[7:0] dcache_io_cpu_resp_bits_tag;
  wire[3:0] dcache_io_cpu_resp_bits_cmd;
  wire[43:0] dcache_io_cpu_resp_bits_addr;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[7:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ptw_req_valid;
  wire[29:0] dcache_io_cpu_ptw_req_bits;
  wire dcache_io_cpu_ordered;
  wire dcache_io_mem_acquire_valid;
  wire[1:0] dcache_io_mem_acquire_bits_header_src;
  wire[1:0] dcache_io_mem_acquire_bits_header_dst;
  wire[25:0] dcache_io_mem_acquire_bits_payload_addr;
  wire[1:0] dcache_io_mem_acquire_bits_payload_client_xact_id;
  wire[135:0] dcache_io_mem_acquire_bits_payload_data;
  wire dcache_io_mem_acquire_bits_payload_uncached;
  wire[1:0] dcache_io_mem_acquire_bits_payload_a_type;
  wire[128:0] dcache_io_mem_acquire_bits_payload_subblock;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_finish_valid;
  wire[1:0] dcache_io_mem_finish_bits_header_src;
  wire[1:0] dcache_io_mem_finish_bits_header_dst;
  wire[3:0] dcache_io_mem_finish_bits_payload_manager_xact_id;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_header_src;
  wire[1:0] dcache_io_mem_release_bits_header_dst;
  wire[25:0] dcache_io_mem_release_bits_payload_addr;
  wire[1:0] dcache_io_mem_release_bits_payload_client_xact_id;
  wire[135:0] dcache_io_mem_release_bits_payload_data;
  wire[2:0] dcache_io_mem_release_bits_payload_r_type;
  wire core_io_host_pcr_req_ready;
  wire core_io_host_pcr_rep_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_pcr;
  wire core_io_imem_req_valid;
  wire[43:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_bits_mask;
  wire core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire[42:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[42:0] core_io_imem_btb_update_bits_pc;
  wire[42:0] core_io_imem_btb_update_bits_target;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isReturn;
  wire[42:0] core_io_imem_btb_update_bits_br_pc;
  wire core_io_imem_bht_update_valid;
  wire core_io_imem_bht_update_bits_prediction_valid;
  wire core_io_imem_bht_update_bits_prediction_bits_taken;
  wire core_io_imem_bht_update_bits_prediction_bits_mask;
  wire core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire[42:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire[42:0] core_io_imem_bht_update_bits_pc;
  wire core_io_imem_bht_update_bits_taken;
  wire core_io_imem_bht_update_bits_mispredict;
  wire core_io_imem_ras_update_valid;
  wire core_io_imem_ras_update_bits_isCall;
  wire core_io_imem_ras_update_bits_isReturn;
  wire[42:0] core_io_imem_ras_update_bits_returnAddr;
  wire core_io_imem_ras_update_bits_prediction_valid;
  wire core_io_imem_ras_update_bits_prediction_bits_taken;
  wire core_io_imem_ras_update_bits_prediction_bits_mask;
  wire core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire[42:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire[5:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire[6:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire core_io_dmem_req_bits_kill;
  wire[3:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_phys;
  wire[43:0] core_io_dmem_req_bits_addr;
  wire[7:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[63:0] core_io_dmem_req_bits_data;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_sret;
  wire[7:0] core_io_ptw_status_ip;
  wire[7:0] core_io_ptw_status_im;
  wire[6:0] core_io_ptw_status_zero;
  wire core_io_ptw_status_er;
  wire core_io_ptw_status_vm;
  wire core_io_ptw_status_s64;
  wire core_io_ptw_status_u64;
  wire core_io_ptw_status_ef;
  wire core_io_ptw_status_pei;
  wire core_io_ptw_status_ei;
  wire core_io_ptw_status_ps;
  wire core_io_ptw_status_s;


  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_tilelink_release_bits_payload_r_type = memArb_io_out_release_bits_payload_r_type;
  assign io_tilelink_release_bits_payload_data = memArb_io_out_release_bits_payload_data;
  assign io_tilelink_release_bits_payload_client_xact_id = memArb_io_out_release_bits_payload_client_xact_id;
  assign io_tilelink_release_bits_payload_addr = memArb_io_out_release_bits_payload_addr;
  assign io_tilelink_release_bits_header_dst = memArb_io_out_release_bits_header_dst;
  assign io_tilelink_release_bits_header_src = memArb_io_out_release_bits_header_src;
  assign io_tilelink_release_valid = memArb_io_out_release_valid;
  assign io_tilelink_probe_ready = memArb_io_out_probe_ready;
  assign io_tilelink_finish_bits_payload_manager_xact_id = memArb_io_out_finish_bits_payload_manager_xact_id;
  assign io_tilelink_finish_bits_header_dst = memArb_io_out_finish_bits_header_dst;
  assign io_tilelink_finish_bits_header_src = memArb_io_out_finish_bits_header_src;
  assign io_tilelink_finish_valid = memArb_io_out_finish_valid;
  assign io_tilelink_grant_ready = memArb_io_out_grant_ready;
  assign io_tilelink_acquire_bits_payload_subblock = memArb_io_out_acquire_bits_payload_subblock;
  assign io_tilelink_acquire_bits_payload_a_type = memArb_io_out_acquire_bits_payload_a_type;
  assign io_tilelink_acquire_bits_payload_uncached = memArb_io_out_acquire_bits_payload_uncached;
  assign io_tilelink_acquire_bits_payload_data = memArb_io_out_acquire_bits_payload_data;
  assign io_tilelink_acquire_bits_payload_client_xact_id = memArb_io_out_acquire_bits_payload_client_xact_id;
  assign io_tilelink_acquire_bits_payload_addr = memArb_io_out_acquire_bits_payload_addr;
  assign io_tilelink_acquire_bits_header_dst = memArb_io_out_acquire_bits_header_dst;
  assign io_tilelink_acquire_bits_header_src = memArb_io_out_acquire_bits_header_src;
  assign io_tilelink_acquire_valid = memArb_io_out_acquire_valid;
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_cpu_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_cpu_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_cpu_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_cpu_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_cpu_btb_update_bits_taken(  )
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_cpu_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_cpu_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_cpu_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_cpu_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_cpu_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_cpu_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_cpu_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_cpu_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_cpu_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_cpu_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_cpu_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_cpu_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_cpu_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_cpu_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_cpu_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_cpu_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_cpu_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_cpu_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_cpu_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_cpu_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_cpu_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_cpu_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_cpu_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_cpu_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_cpu_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_0_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_0_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_0_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_0_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_0_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_0_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_0_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_0_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_0_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_0_sret ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_mem_acquire_ready( TileLinkIOWrapper_io_in_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( icache_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( icache_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( TileLinkIOWrapper_io_in_grant_valid ),
       .io_mem_grant_bits_header_src( TileLinkIOWrapper_io_in_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( TileLinkIOWrapper_io_in_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( TileLinkIOWrapper_io_in_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( TileLinkIOWrapper_io_in_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( TileLinkIOWrapper_io_in_grant_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( TileLinkIOWrapper_io_in_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( TileLinkIOWrapper_io_in_grant_bits_payload_g_type ),
       .io_mem_finish_ready( TileLinkIOWrapper_io_in_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( icache_io_mem_finish_bits_payload_manager_xact_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign icache.io_cpu_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_cpu_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_1_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_1_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_1_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_1_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_1_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_1_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_1_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_1_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_1_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_1_sret ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_mem_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_mem_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_mem_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( dcache_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( dcache_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_0_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( memArb_io_in_0_grant_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( memArb_io_in_0_grant_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_0_finish_ready ),
       .io_mem_finish_valid( dcache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( dcache_io_mem_finish_bits_payload_manager_xact_id ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( memArb_io_in_0_probe_valid ),
       .io_mem_probe_bits_header_src( memArb_io_in_0_probe_bits_header_src ),
       .io_mem_probe_bits_header_dst( memArb_io_in_0_probe_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( memArb_io_in_0_probe_bits_payload_addr ),
       .io_mem_probe_bits_payload_p_type( memArb_io_in_0_probe_bits_payload_p_type ),
       .io_mem_release_ready( memArb_io_in_0_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_mem_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_mem_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_requestor_1_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_requestor_1_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_requestor_1_status_ip( ptw_io_requestor_1_status_ip ),
       .io_requestor_1_status_im( ptw_io_requestor_1_status_im ),
       .io_requestor_1_status_zero( ptw_io_requestor_1_status_zero ),
       .io_requestor_1_status_er( ptw_io_requestor_1_status_er ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_requestor_1_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_requestor_1_status_ef( ptw_io_requestor_1_status_ef ),
       .io_requestor_1_status_pei( ptw_io_requestor_1_status_pei ),
       .io_requestor_1_status_ei( ptw_io_requestor_1_status_ei ),
       .io_requestor_1_status_ps( ptw_io_requestor_1_status_ps ),
       .io_requestor_1_status_s( ptw_io_requestor_1_status_s ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_1_sret( ptw_io_requestor_1_sret ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_requestor_0_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_requestor_0_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_requestor_0_status_ip( ptw_io_requestor_0_status_ip ),
       .io_requestor_0_status_im( ptw_io_requestor_0_status_im ),
       .io_requestor_0_status_zero( ptw_io_requestor_0_status_zero ),
       .io_requestor_0_status_er( ptw_io_requestor_0_status_er ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_requestor_0_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_requestor_0_status_ef( ptw_io_requestor_0_status_ef ),
       .io_requestor_0_status_pei( ptw_io_requestor_0_status_pei ),
       .io_requestor_0_status_ei( ptw_io_requestor_0_status_ei ),
       .io_requestor_0_status_ps( ptw_io_requestor_0_status_ps ),
       .io_requestor_0_status_s( ptw_io_requestor_0_status_s ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_requestor_0_sret( ptw_io_requestor_0_sret ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       //.io_mem_req_bits_data(  )
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       //.io_mem_ptw_req_valid(  )
       //.io_mem_ptw_req_bits(  )
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_sret( core_io_ptw_sret ),
       .io_dpath_status_ip( core_io_ptw_status_ip ),
       .io_dpath_status_im( core_io_ptw_status_im ),
       .io_dpath_status_zero( core_io_ptw_status_zero ),
       .io_dpath_status_er( core_io_ptw_status_er ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_s64( core_io_ptw_status_s64 ),
       .io_dpath_status_u64( core_io_ptw_status_u64 ),
       .io_dpath_status_ef( core_io_ptw_status_ef ),
       .io_dpath_status_pei( core_io_ptw_status_pei ),
       .io_dpath_status_ei( core_io_ptw_status_ei ),
       .io_dpath_status_ps( core_io_ptw_status_ps ),
       .io_dpath_status_s( core_io_ptw_status_s )
  );
  Core core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_imem_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_imem_btb_update_bits_taken(  )
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_imem_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_imem_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_imem_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_imem_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_imem_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_imem_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_imem_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_imem_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_imem_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_imem_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_imem_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_imem_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_imem_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_imem_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_imem_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_imem_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_imem_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_imem_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_imem_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_imem_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_imem_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_imem_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_imem_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_imem_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_imem_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       //.io_dmem_ptw_req_valid(  )
       //.io_dmem_ptw_req_bits(  )
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_sret( core_io_ptw_sret ),
       .io_ptw_status_ip( core_io_ptw_status_ip ),
       .io_ptw_status_im( core_io_ptw_status_im ),
       .io_ptw_status_zero( core_io_ptw_status_zero ),
       .io_ptw_status_er( core_io_ptw_status_er ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_s64( core_io_ptw_status_s64 ),
       .io_ptw_status_u64( core_io_ptw_status_u64 ),
       .io_ptw_status_ef( core_io_ptw_status_ef ),
       .io_ptw_status_pei( core_io_ptw_status_pei ),
       .io_ptw_status_ei( core_io_ptw_status_ei ),
       .io_ptw_status_ps( core_io_ptw_status_ps ),
       .io_ptw_status_s( core_io_ptw_status_s )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_uncached(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_subblock(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_uncached(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       //.io_rocc_imem_finish_valid(  )
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_manager_xact_id(  )
       //.io_rocc_dmem_acquire_ready(  )
       //.io_rocc_dmem_acquire_valid(  )
       //.io_rocc_dmem_acquire_bits_header_src(  )
       //.io_rocc_dmem_acquire_bits_header_dst(  )
       //.io_rocc_dmem_acquire_bits_payload_addr(  )
       //.io_rocc_dmem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_dmem_acquire_bits_payload_data(  )
       //.io_rocc_dmem_acquire_bits_payload_uncached(  )
       //.io_rocc_dmem_acquire_bits_payload_a_type(  )
       //.io_rocc_dmem_acquire_bits_payload_subblock(  )
       //.io_rocc_dmem_grant_ready(  )
       //.io_rocc_dmem_grant_valid(  )
       //.io_rocc_dmem_grant_bits_header_src(  )
       //.io_rocc_dmem_grant_bits_header_dst(  )
       //.io_rocc_dmem_grant_bits_payload_data(  )
       //.io_rocc_dmem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_manager_xact_id(  )
       //.io_rocc_dmem_grant_bits_payload_uncached(  )
       //.io_rocc_dmem_grant_bits_payload_g_type(  )
       //.io_rocc_dmem_finish_ready(  )
       //.io_rocc_dmem_finish_valid(  )
       //.io_rocc_dmem_finish_bits_header_src(  )
       //.io_rocc_dmem_finish_bits_header_dst(  )
       //.io_rocc_dmem_finish_bits_payload_manager_xact_id(  )
       //.io_rocc_dmem_probe_ready(  )
       //.io_rocc_dmem_probe_valid(  )
       //.io_rocc_dmem_probe_bits_header_src(  )
       //.io_rocc_dmem_probe_bits_header_dst(  )
       //.io_rocc_dmem_probe_bits_payload_addr(  )
       //.io_rocc_dmem_probe_bits_payload_p_type(  )
       //.io_rocc_dmem_release_ready(  )
       //.io_rocc_dmem_release_valid(  )
       //.io_rocc_dmem_release_bits_header_src(  )
       //.io_rocc_dmem_release_bits_header_dst(  )
       //.io_rocc_dmem_release_bits_payload_addr(  )
       //.io_rocc_dmem_release_bits_payload_client_xact_id(  )
       //.io_rocc_dmem_release_bits_payload_data(  )
       //.io_rocc_dmem_release_bits_payload_r_type(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign core.io_dmem_ptw_req_valid = {1{$random}};
    assign core.io_dmem_ptw_req_bits = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_ptw_req_ready = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_valid = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_error = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_ppn = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_perm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ip = {1{$random}};
    assign core.io_rocc_mem_ptw_status_im = {1{$random}};
    assign core.io_rocc_mem_ptw_status_zero = {1{$random}};
    assign core.io_rocc_mem_ptw_status_er = {1{$random}};
    assign core.io_rocc_mem_ptw_status_vm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_u64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ef = {1{$random}};
    assign core.io_rocc_mem_ptw_status_pei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ps = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s = {1{$random}};
    assign core.io_rocc_mem_ptw_invalidate = {1{$random}};
    assign core.io_rocc_mem_ptw_sret = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_data = {5{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_uncached = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_subblock = {5{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_imem_finish_valid = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_finish_bits_payload_manager_xact_id = {1{$random}};
    assign core.io_rocc_dmem_acquire_valid = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_payload_data = {5{$random}};
    assign core.io_rocc_dmem_acquire_bits_payload_uncached = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_payload_subblock = {5{$random}};
    assign core.io_rocc_dmem_grant_ready = {1{$random}};
    assign core.io_rocc_dmem_finish_valid = {1{$random}};
    assign core.io_rocc_dmem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_dmem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_dmem_finish_bits_payload_manager_xact_id = {1{$random}};
    assign core.io_rocc_dmem_probe_ready = {1{$random}};
    assign core.io_rocc_dmem_release_valid = {1{$random}};
    assign core.io_rocc_dmem_release_bits_header_src = {1{$random}};
    assign core.io_rocc_dmem_release_bits_header_dst = {1{$random}};
    assign core.io_rocc_dmem_release_bits_payload_addr = {1{$random}};
    assign core.io_rocc_dmem_release_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_dmem_release_bits_payload_data = {5{$random}};
    assign core.io_rocc_dmem_release_bits_payload_r_type = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits = {1{$random}};
// synthesis translate_on
`endif
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_requestor_1_ptw_req_ready(  )
       //.io_requestor_1_ptw_req_valid(  )
       //.io_requestor_1_ptw_req_bits(  )
       //.io_requestor_1_ptw_resp_valid(  )
       //.io_requestor_1_ptw_resp_bits_error(  )
       //.io_requestor_1_ptw_resp_bits_ppn(  )
       //.io_requestor_1_ptw_resp_bits_perm(  )
       //.io_requestor_1_ptw_status_ip(  )
       //.io_requestor_1_ptw_status_im(  )
       //.io_requestor_1_ptw_status_zero(  )
       //.io_requestor_1_ptw_status_er(  )
       //.io_requestor_1_ptw_status_vm(  )
       //.io_requestor_1_ptw_status_s64(  )
       //.io_requestor_1_ptw_status_u64(  )
       //.io_requestor_1_ptw_status_ef(  )
       //.io_requestor_1_ptw_status_pei(  )
       //.io_requestor_1_ptw_status_ei(  )
       //.io_requestor_1_ptw_status_ps(  )
       //.io_requestor_1_ptw_status_s(  )
       //.io_requestor_1_ptw_invalidate(  )
       //.io_requestor_1_ptw_sret(  )
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       //.io_requestor_0_req_bits_data(  )
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_ptw_req_ready(  )
       //.io_requestor_0_ptw_req_valid(  )
       //.io_requestor_0_ptw_req_bits(  )
       //.io_requestor_0_ptw_resp_valid(  )
       //.io_requestor_0_ptw_resp_bits_error(  )
       //.io_requestor_0_ptw_resp_bits_ppn(  )
       //.io_requestor_0_ptw_resp_bits_perm(  )
       //.io_requestor_0_ptw_status_ip(  )
       //.io_requestor_0_ptw_status_im(  )
       //.io_requestor_0_ptw_status_zero(  )
       //.io_requestor_0_ptw_status_er(  )
       //.io_requestor_0_ptw_status_vm(  )
       //.io_requestor_0_ptw_status_s64(  )
       //.io_requestor_0_ptw_status_u64(  )
       //.io_requestor_0_ptw_status_ef(  )
       //.io_requestor_0_ptw_status_pei(  )
       //.io_requestor_0_ptw_status_ei(  )
       //.io_requestor_0_ptw_status_ps(  )
       //.io_requestor_0_ptw_status_s(  )
       //.io_requestor_0_ptw_invalidate(  )
       //.io_requestor_0_ptw_sret(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_mem_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
    assign dcArb.io_requestor_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  TileLinkIOArbiterThatAppendsArbiterId memArb(.clk(clk), .reset(reset),
       .io_in_1_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( TileLinkIOWrapper_io_out_acquire_valid ),
       .io_in_1_acquire_bits_header_src( TileLinkIOWrapper_io_out_acquire_bits_header_src ),
       .io_in_1_acquire_bits_header_dst( TileLinkIOWrapper_io_out_acquire_bits_header_dst ),
       .io_in_1_acquire_bits_payload_addr( TileLinkIOWrapper_io_out_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( TileLinkIOWrapper_io_out_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( TileLinkIOWrapper_io_out_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_uncached( TileLinkIOWrapper_io_out_acquire_bits_payload_uncached ),
       .io_in_1_acquire_bits_payload_a_type( TileLinkIOWrapper_io_out_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_subblock( TileLinkIOWrapper_io_out_acquire_bits_payload_subblock ),
       .io_in_1_grant_ready( TileLinkIOWrapper_io_out_grant_ready ),
       .io_in_1_grant_valid( memArb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_manager_xact_id( memArb_io_in_1_grant_bits_payload_manager_xact_id ),
       .io_in_1_grant_bits_payload_uncached( memArb_io_in_1_grant_bits_payload_uncached ),
       .io_in_1_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( memArb_io_in_1_finish_ready ),
       .io_in_1_finish_valid( TileLinkIOWrapper_io_out_finish_valid ),
       .io_in_1_finish_bits_header_src( TileLinkIOWrapper_io_out_finish_bits_header_src ),
       .io_in_1_finish_bits_header_dst( TileLinkIOWrapper_io_out_finish_bits_header_dst ),
       .io_in_1_finish_bits_payload_manager_xact_id( TileLinkIOWrapper_io_out_finish_bits_payload_manager_xact_id ),
       .io_in_1_probe_ready( TileLinkIOWrapper_io_out_probe_ready ),
       .io_in_1_probe_valid( memArb_io_in_1_probe_valid ),
       .io_in_1_probe_bits_header_src( memArb_io_in_1_probe_bits_header_src ),
       .io_in_1_probe_bits_header_dst( memArb_io_in_1_probe_bits_header_dst ),
       .io_in_1_probe_bits_payload_addr( memArb_io_in_1_probe_bits_payload_addr ),
       .io_in_1_probe_bits_payload_p_type( memArb_io_in_1_probe_bits_payload_p_type ),
       .io_in_1_release_ready( memArb_io_in_1_release_ready ),
       .io_in_1_release_valid( TileLinkIOWrapper_io_out_release_valid ),
       //.io_in_1_release_bits_header_src(  )
       //.io_in_1_release_bits_header_dst(  )
       //.io_in_1_release_bits_payload_addr(  )
       //.io_in_1_release_bits_payload_client_xact_id(  )
       //.io_in_1_release_bits_payload_data(  )
       //.io_in_1_release_bits_payload_r_type(  )
       .io_in_0_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_in_0_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_in_0_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_uncached( dcache_io_mem_acquire_bits_payload_uncached ),
       .io_in_0_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_subblock( dcache_io_mem_acquire_bits_payload_subblock ),
       .io_in_0_grant_ready( dcache_io_mem_grant_ready ),
       .io_in_0_grant_valid( memArb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_manager_xact_id( memArb_io_in_0_grant_bits_payload_manager_xact_id ),
       .io_in_0_grant_bits_payload_uncached( memArb_io_in_0_grant_bits_payload_uncached ),
       .io_in_0_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( memArb_io_in_0_finish_ready ),
       .io_in_0_finish_valid( dcache_io_mem_finish_valid ),
       .io_in_0_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_in_0_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_in_0_finish_bits_payload_manager_xact_id( dcache_io_mem_finish_bits_payload_manager_xact_id ),
       .io_in_0_probe_ready( dcache_io_mem_probe_ready ),
       .io_in_0_probe_valid( memArb_io_in_0_probe_valid ),
       .io_in_0_probe_bits_header_src( memArb_io_in_0_probe_bits_header_src ),
       .io_in_0_probe_bits_header_dst( memArb_io_in_0_probe_bits_header_dst ),
       .io_in_0_probe_bits_payload_addr( memArb_io_in_0_probe_bits_payload_addr ),
       .io_in_0_probe_bits_payload_p_type( memArb_io_in_0_probe_bits_payload_p_type ),
       .io_in_0_release_ready( memArb_io_in_0_release_ready ),
       .io_in_0_release_valid( dcache_io_mem_release_valid ),
       .io_in_0_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_in_0_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_in_0_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_in_0_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_in_0_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_in_0_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type ),
       .io_out_acquire_ready( io_tilelink_acquire_ready ),
       .io_out_acquire_valid( memArb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( memArb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( memArb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( memArb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( memArb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( memArb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_uncached( memArb_io_out_acquire_bits_payload_uncached ),
       .io_out_acquire_bits_payload_a_type( memArb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_subblock( memArb_io_out_acquire_bits_payload_subblock ),
       .io_out_grant_ready( memArb_io_out_grant_ready ),
       .io_out_grant_valid( io_tilelink_grant_valid ),
       .io_out_grant_bits_header_src( io_tilelink_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_tilelink_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_tilelink_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_tilelink_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_manager_xact_id( io_tilelink_grant_bits_payload_manager_xact_id ),
       .io_out_grant_bits_payload_uncached( io_tilelink_grant_bits_payload_uncached ),
       .io_out_grant_bits_payload_g_type( io_tilelink_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_tilelink_finish_ready ),
       .io_out_finish_valid( memArb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( memArb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( memArb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_manager_xact_id( memArb_io_out_finish_bits_payload_manager_xact_id ),
       .io_out_probe_ready( memArb_io_out_probe_ready ),
       .io_out_probe_valid( io_tilelink_probe_valid ),
       .io_out_probe_bits_header_src( io_tilelink_probe_bits_header_src ),
       .io_out_probe_bits_header_dst( io_tilelink_probe_bits_header_dst ),
       .io_out_probe_bits_payload_addr( io_tilelink_probe_bits_payload_addr ),
       .io_out_probe_bits_payload_p_type( io_tilelink_probe_bits_payload_p_type ),
       .io_out_release_ready( io_tilelink_release_ready ),
       .io_out_release_valid( memArb_io_out_release_valid ),
       .io_out_release_bits_header_src( memArb_io_out_release_bits_header_src ),
       .io_out_release_bits_header_dst( memArb_io_out_release_bits_header_dst ),
       .io_out_release_bits_payload_addr( memArb_io_out_release_bits_payload_addr ),
       .io_out_release_bits_payload_client_xact_id( memArb_io_out_release_bits_payload_client_xact_id ),
       .io_out_release_bits_payload_data( memArb_io_out_release_bits_payload_data ),
       .io_out_release_bits_payload_r_type( memArb_io_out_release_bits_payload_r_type )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign memArb.io_in_1_release_bits_header_src = {1{$random}};
    assign memArb.io_in_1_release_bits_header_dst = {1{$random}};
    assign memArb.io_in_1_release_bits_payload_addr = {1{$random}};
    assign memArb.io_in_1_release_bits_payload_client_xact_id = {1{$random}};
    assign memArb.io_in_1_release_bits_payload_data = {5{$random}};
    assign memArb.io_in_1_release_bits_payload_r_type = {1{$random}};
// synthesis translate_on
`endif
  TileLinkIOWrapper TileLinkIOWrapper(
       .io_in_acquire_ready( TileLinkIOWrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_in_acquire_bits_header_src(  )
       //.io_in_acquire_bits_header_dst(  )
       .io_in_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_in_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_in_acquire_bits_payload_uncached( icache_io_mem_acquire_bits_payload_uncached ),
       .io_in_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_in_acquire_bits_payload_subblock( icache_io_mem_acquire_bits_payload_subblock ),
       .io_in_grant_ready( icache_io_mem_grant_ready ),
       .io_in_grant_valid( TileLinkIOWrapper_io_in_grant_valid ),
       .io_in_grant_bits_header_src( TileLinkIOWrapper_io_in_grant_bits_header_src ),
       .io_in_grant_bits_header_dst( TileLinkIOWrapper_io_in_grant_bits_header_dst ),
       .io_in_grant_bits_payload_data( TileLinkIOWrapper_io_in_grant_bits_payload_data ),
       .io_in_grant_bits_payload_client_xact_id( TileLinkIOWrapper_io_in_grant_bits_payload_client_xact_id ),
       .io_in_grant_bits_payload_manager_xact_id( TileLinkIOWrapper_io_in_grant_bits_payload_manager_xact_id ),
       .io_in_grant_bits_payload_uncached( TileLinkIOWrapper_io_in_grant_bits_payload_uncached ),
       .io_in_grant_bits_payload_g_type( TileLinkIOWrapper_io_in_grant_bits_payload_g_type ),
       .io_in_finish_ready( TileLinkIOWrapper_io_in_finish_ready ),
       .io_in_finish_valid( icache_io_mem_finish_valid ),
       .io_in_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_in_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_in_finish_bits_payload_manager_xact_id( icache_io_mem_finish_bits_payload_manager_xact_id ),
       .io_out_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_out_acquire_valid( TileLinkIOWrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( TileLinkIOWrapper_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( TileLinkIOWrapper_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( TileLinkIOWrapper_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( TileLinkIOWrapper_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( TileLinkIOWrapper_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_uncached( TileLinkIOWrapper_io_out_acquire_bits_payload_uncached ),
       .io_out_acquire_bits_payload_a_type( TileLinkIOWrapper_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_subblock( TileLinkIOWrapper_io_out_acquire_bits_payload_subblock ),
       .io_out_grant_ready( TileLinkIOWrapper_io_out_grant_ready ),
       .io_out_grant_valid( memArb_io_in_1_grant_valid ),
       .io_out_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_manager_xact_id( memArb_io_in_1_grant_bits_payload_manager_xact_id ),
       .io_out_grant_bits_payload_uncached( memArb_io_in_1_grant_bits_payload_uncached ),
       .io_out_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_out_finish_ready( memArb_io_in_1_finish_ready ),
       .io_out_finish_valid( TileLinkIOWrapper_io_out_finish_valid ),
       .io_out_finish_bits_header_src( TileLinkIOWrapper_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( TileLinkIOWrapper_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_manager_xact_id( TileLinkIOWrapper_io_out_finish_bits_payload_manager_xact_id ),
       .io_out_probe_ready( TileLinkIOWrapper_io_out_probe_ready ),
       .io_out_probe_valid( memArb_io_in_1_probe_valid ),
       .io_out_probe_bits_header_src( memArb_io_in_1_probe_bits_header_src ),
       .io_out_probe_bits_header_dst( memArb_io_in_1_probe_bits_header_dst ),
       .io_out_probe_bits_payload_addr( memArb_io_in_1_probe_bits_payload_addr ),
       .io_out_probe_bits_payload_p_type( memArb_io_in_1_probe_bits_payload_p_type ),
       .io_out_release_ready( memArb_io_in_1_release_ready ),
       .io_out_release_valid( TileLinkIOWrapper_io_out_release_valid )
       //.io_out_release_bits_header_src(  )
       //.io_out_release_bits_header_dst(  )
       //.io_out_release_bits_payload_addr(  )
       //.io_out_release_bits_payload_client_xact_id(  )
       //.io_out_release_bits_payload_data(  )
       //.io_out_release_bits_payload_r_type(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign TileLinkIOWrapper.io_in_acquire_bits_header_src = {1{$random}};
    assign TileLinkIOWrapper.io_in_acquire_bits_header_dst = {1{$random}};
// synthesis translate_on
`endif
endmodule

module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[4:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[135:0] io_mem_acquire_bits_payload_data,
    output io_mem_acquire_bits_payload_uncached,
    output[1:0] io_mem_acquire_bits_payload_a_type,
    output[128:0] io_mem_acquire_bits_payload_subblock,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [135:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_manager_xact_id,
    input  io_mem_grant_bits_payload_uncached,
    input [1:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    //output[1:0] io_mem_finish_bits_header_src
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_manager_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    //output[1:0] io_mem_release_bits_header_src
    //output[1:0] io_mem_release_bits_header_dst
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[135:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[63:0] pcr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire[127:0] grant_payload_without_tag;
  wire[127:0] T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire T5;
  wire T6;
  reg [3:0] state;
  wire[3:0] T340;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire[3:0] rx_cmd;
  reg [3:0] cmd;
  wire[3:0] T23;
  wire T24;
  wire T25;
  reg [14:0] rx_count;
  wire[14:0] T341;
  wire[14:0] T26;
  wire[14:0] T27;
  wire[14:0] T28;
  wire T29;
  wire T30;
  wire[12:0] T342;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T31;
  wire[11:0] T32;
  wire[63:0] rx_shifter_in;
  wire[47:0] T33;
  reg [63:0] rx_shifter;
  wire[63:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire nack;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire bad_mem_packet;
  wire T47;
  wire[2:0] T48;
  reg [39:0] addr;
  wire[39:0] T49;
  wire[39:0] T50;
  wire[39:0] T51;
  wire[39:0] T52;
  wire T53;
  wire[2:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T343;
  wire[14:0] T58;
  wire[14:0] T59;
  wire[14:0] T60;
  wire T61;
  wire T62;
  wire[3:0] next_cmd;
  wire T63;
  wire[12:0] rx_word_count;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire rx_done;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire T72;
  wire[12:0] T344;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire rx_word_done;
  wire T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire cnt_done;
  wire T81;
  reg [1:0] cnt;
  wire[1:0] T345;
  wire[1:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg  mem_acked;
  wire T346;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[3:0] T99;
  wire T100;
  wire T101;
  reg [8:0] pos;
  wire[8:0] T102;
  wire[8:0] T103;
  wire[8:0] T104;
  wire[8:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire[3:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire tx_done;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire[12:0] T347;
  wire T120;
  wire T121;
  wire[1:0] tx_subword_count;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[4:0] pcr_addr;
  wire T126;
  wire T127;
  wire[1:0] pcr_coreid;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire[63:0] T133;
  wire[63:0] T134;
  wire T135;
  wire T136;
  wire[2:0] T137;
  wire[63:0] T138;
  wire T139;
  wire[2:0] T140;
  wire[2:0] T141;
  wire[5:0] T142;
  wire[5:0] scr_addr;
  wire T143;
  wire T144;
  reg [3:0] mem_gxid;
  wire[3:0] T145;
  reg [1:0] mem_gsrc;
  wire[1:0] T146;
  wire T147;
  reg  mem_needs_ack;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[128:0] T152;
  wire[128:0] T153;
  wire[128:0] T154;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire[135:0] T162;
  wire[135:0] T163;
  wire[67:0] T164;
  wire[63:0] T165;
  wire[127:0] mem_req_data;
  wire[63:0] T166;
  wire[63:0] T167;
  wire[67:0] T168;
  wire[63:0] T169;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire[25:0] T173;
  wire[25:0] T174;
  wire[25:0] T348;
  wire[36:0] init_addr;
  wire[39:0] T175;
  wire[25:0] T176;
  wire[25:0] T349;
  wire T177;
  wire T178;
  wire T179;
  reg  R180;
  wire T350;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  reg  R190;
  wire T351;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire[15:0] T352;
  wire[63:0] T195;
  wire[5:0] T196;
  wire[1:0] T197;
  wire[63:0] tx_data;
  wire[63:0] T198;
  wire[63:0] T199;
  reg [63:0] pcrReadData;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  wire[63:0] T353;
  wire[63:0] T203;
  wire[63:0] T204;
  wire[63:0] T205;
  wire[63:0] T206;
  wire[63:0] T207;
  wire[63:0] T208;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T209;
  wire[5:0] T210;
  wire[63:0] T211;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T212;
  wire T213;
  wire[63:0] T214;
  wire[63:0] T215;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T216;
  wire[63:0] T217;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T218;
  wire T219;
  wire T220;
  wire[63:0] T221;
  wire[63:0] T222;
  wire[63:0] T223;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T224;
  wire[63:0] T225;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T226;
  wire T227;
  wire[63:0] T228;
  wire[63:0] T229;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T230;
  wire[63:0] T231;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire[63:0] T236;
  wire[63:0] T237;
  wire[63:0] T238;
  wire[63:0] T239;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T240;
  wire[63:0] T241;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T242;
  wire T243;
  wire[63:0] T244;
  wire[63:0] T245;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T246;
  wire[63:0] T247;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T248;
  wire T249;
  wire T250;
  wire[63:0] T251;
  wire[63:0] T252;
  wire[63:0] T253;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T254;
  wire[63:0] T255;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T256;
  wire T257;
  wire[63:0] T258;
  wire[63:0] T259;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T260;
  wire[63:0] T261;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire[63:0] T267;
  wire[63:0] T268;
  wire[63:0] T269;
  wire[63:0] T270;
  wire[63:0] T271;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T272;
  wire[63:0] T273;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T274;
  wire T275;
  wire[63:0] T276;
  wire[63:0] T277;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T278;
  wire[63:0] T279;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T280;
  wire T281;
  wire T282;
  wire[63:0] T283;
  wire[63:0] T284;
  wire[63:0] T285;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T286;
  wire[63:0] T287;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T288;
  wire T289;
  wire[63:0] T290;
  wire[63:0] T291;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T292;
  wire[63:0] T293;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[63:0] T298;
  wire[63:0] T299;
  wire[63:0] T300;
  wire[63:0] T301;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T302;
  wire[63:0] T303;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T304;
  wire T305;
  wire[63:0] T306;
  wire[63:0] T307;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T308;
  wire[63:0] T309;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T310;
  wire T311;
  wire T312;
  wire[63:0] T313;
  wire[63:0] T314;
  wire[63:0] T315;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T316;
  wire[63:0] T317;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T318;
  wire T319;
  wire[63:0] T320;
  wire[63:0] T321;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T322;
  wire[63:0] T323;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire[63:0] tx_header;
  wire[15:0] T333;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T334;
  reg [7:0] seqno;
  wire[7:0] T335;
  wire[7:0] T336;
  wire T337;
  wire T338;
  wire T339;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    state = {1{$random}};
    cmd = {1{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    rx_shifter = {2{$random}};
    addr = {2{$random}};
    tx_count = {1{$random}};
    cnt = {1{$random}};
    mem_acked = {1{$random}};
    pos = {1{$random}};
    mem_gxid = {1{$random}};
    mem_gsrc = {1{$random}};
    mem_needs_ack = {1{$random}};
    R180 = {1{$random}};
    R190 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_scr_wdata = pcr_wdata;
  assign pcr_wdata = packet_ram[3'h0];
  assign T1 = grant_payload_without_tag[7'h7f:7'h40];
  assign grant_payload_without_tag = T2;
  assign T2 = {T4, T3};
  assign T3 = io_mem_grant_bits_payload_data[6'h3f:1'h0];
  assign T4 = io_mem_grant_bits_payload_data[8'h83:7'h44];
  assign T5 = T6 & io_mem_grant_valid;
  assign T6 = state == 4'h5;
  assign T340 = reset ? 4'h0 : T7;
  assign T7 = T129 ? 4'h8 : T8;
  assign T8 = io_cpu_0_pcr_rep_valid ? 4'h8 : T9;
  assign T9 = T124 ? 4'h8 : T10;
  assign T10 = T123 ? 4'h2 : T11;
  assign T11 = T113 ? T109 : T12;
  assign T12 = T107 ? T99 : T13;
  assign T13 = T97 ? 4'h7 : T14;
  assign T14 = T92 ? 4'h7 : T15;
  assign T15 = T90 ? 4'h5 : T16;
  assign T16 = T80 ? 4'h6 : T17;
  assign T17 = T67 ? T18 : state;
  assign T18 = T66 ? 4'h3 : T19;
  assign T19 = T65 ? 4'h4 : T20;
  assign T20 = T21 ? 4'h1 : 4'h8;
  assign T21 = T64 | T22;
  assign T22 = rx_cmd == 4'h3;
  assign rx_cmd = T63 ? next_cmd : cmd;
  assign T23 = T24 ? next_cmd : cmd;
  assign T24 = T62 & T25;
  assign T25 = rx_count == 15'h3;
  assign T341 = reset ? 15'h0 : T26;
  assign T26 = T29 ? 15'h0 : T27;
  assign T27 = T62 ? T28 : rx_count;
  assign T28 = rx_count + 15'h1;
  assign T29 = T113 & T30;
  assign T30 = tx_word_count == T342;
  assign T342 = {1'h0, tx_size};
  assign tx_size = T35 ? size : 12'h0;
  assign T31 = T24 ? T32 : size;
  assign T32 = rx_shifter_in[4'hf:3'h4];
  assign rx_shifter_in = {io_host_in_bits, T33};
  assign T33 = rx_shifter[6'h3f:5'h10];
  assign T34 = T62 ? rx_shifter_in : rx_shifter;
  assign T35 = T41 & T36;
  assign T36 = T38 | T37;
  assign T37 = cmd == 4'h3;
  assign T38 = T40 | T39;
  assign T39 = cmd == 4'h2;
  assign T40 = cmd == 4'h0;
  assign T41 = nack ^ 1'h1;
  assign nack = T55 ? bad_mem_packet : T42;
  assign T42 = T44 ? T43 : 1'h1;
  assign T43 = size != 12'h1;
  assign T44 = T46 | T45;
  assign T45 = cmd == 4'h3;
  assign T46 = cmd == 4'h2;
  assign bad_mem_packet = T53 | T47;
  assign T47 = T48 != 3'h0;
  assign T48 = addr[2'h2:1'h0];
  assign T49 = T107 ? T52 : T50;
  assign T50 = T24 ? T51 : addr;
  assign T51 = rx_shifter_in[6'h3f:5'h18];
  assign T52 = addr + 40'h8;
  assign T53 = T54 != 3'h0;
  assign T54 = size[2'h2:1'h0];
  assign T55 = T57 | T56;
  assign T56 = cmd == 4'h1;
  assign T57 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T343 = reset ? 15'h0 : T58;
  assign T58 = T29 ? 15'h0 : T59;
  assign T59 = T61 ? T60 : tx_count;
  assign T60 = tx_count + 15'h1;
  assign T61 = io_host_out_valid & io_host_out_ready;
  assign T62 = io_host_in_valid & io_host_in_ready;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign T63 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T64 = rx_cmd == 4'h2;
  assign T65 = rx_cmd == 4'h1;
  assign T66 = rx_cmd == 4'h0;
  assign T67 = T79 & rx_done;
  assign rx_done = rx_word_done & T68;
  assign T68 = T76 ? T73 : T69;
  assign T69 = T72 | T70;
  assign T70 = T71 == 3'h0;
  assign T71 = rx_word_count[2'h2:1'h0];
  assign T72 = rx_word_count == T344;
  assign T344 = {1'h0, size};
  assign T73 = T75 & T74;
  assign T74 = next_cmd != 4'h3;
  assign T75 = next_cmd != 4'h1;
  assign T76 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T77;
  assign T77 = T78 == 2'h3;
  assign T78 = rx_count[1'h1:1'h0];
  assign T79 = state == 4'h0;
  assign T80 = T89 & cnt_done;
  assign cnt_done = T84 & T81;
  assign T81 = cnt == 2'h3;
  assign T345 = reset ? 2'h0 : T82;
  assign T82 = T84 ? T83 : cnt;
  assign T83 = cnt + 2'h1;
  assign T84 = T87 | T85;
  assign T85 = T86 & io_mem_grant_valid;
  assign T86 = state == 4'h5;
  assign T87 = T88 & io_mem_acquire_ready;
  assign T88 = state == 4'h4;
  assign T89 = state == 4'h4;
  assign T90 = T91 & io_mem_acquire_ready;
  assign T91 = state == 4'h3;
  assign T92 = T96 & mem_acked;
  assign T346 = reset ? 1'h0 : T93;
  assign T93 = T97 ? 1'h0 : T94;
  assign T94 = T92 ? 1'h0 : T95;
  assign T95 = io_mem_grant_valid ? 1'h1 : mem_acked;
  assign T96 = state == 4'h6;
  assign T97 = T98 & cnt_done;
  assign T98 = state == 4'h5;
  assign T99 = T100 ? 4'h8 : 4'h0;
  assign T100 = T106 | T101;
  assign T101 = pos == 9'h1;
  assign T102 = T107 ? T105 : T103;
  assign T103 = T24 ? T104 : pos;
  assign T104 = rx_shifter_in[4'hf:3'h7];
  assign T105 = pos - 9'h1;
  assign T106 = cmd == 4'h0;
  assign T107 = T108 & io_mem_finish_ready;
  assign T108 = state == 4'h7;
  assign T109 = T110 ? 4'h3 : 4'h0;
  assign T110 = T112 & T111;
  assign T111 = pos != 9'h0;
  assign T112 = cmd == 4'h0;
  assign T113 = T122 & tx_done;
  assign tx_done = T120 & T114;
  assign T114 = T119 | T115;
  assign T115 = T118 & T116;
  assign T116 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T117 - 3'h1;
  assign T117 = tx_word_count[2'h2:1'h0];
  assign T118 = 13'h0 < tx_word_count;
  assign T119 = tx_word_count == T347;
  assign T347 = {1'h0, tx_size};
  assign T120 = io_host_out_ready & T121;
  assign T121 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T122 = state == 4'h8;
  assign T123 = io_cpu_0_pcr_req_valid & io_cpu_0_pcr_req_ready;
  assign T124 = T126 & T125;
  assign T125 = pcr_addr == 5'h1d;
  assign pcr_addr = addr[3'h4:1'h0];
  assign T126 = T128 & T127;
  assign T127 = pcr_coreid == 2'h0;
  assign pcr_coreid = addr[5'h15:5'h14];
  assign T128 = state == 4'h1;
  assign T129 = T131 & T130;
  assign T130 = pcr_coreid == 2'h3;
  assign T131 = state == 4'h1;
  assign T132 = {cnt, 1'h1};
  assign T134 = grant_payload_without_tag[6'h3f:1'h0];
  assign T135 = T136 & io_mem_grant_valid;
  assign T136 = state == 4'h5;
  assign T137 = {cnt, 1'h0};
  assign T139 = rx_word_done & io_host_in_ready;
  assign T140 = T141 - 3'h1;
  assign T141 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T142;
  assign T142 = scr_addr;
  assign scr_addr = addr[3'h5:1'h0];
  assign io_scr_wen = T143;
  assign T143 = T129 ? T144 : 1'h0;
  assign T144 = cmd == 4'h3;
  assign io_mem_release_bits_payload_r_type = {1{$random}};
  assign io_mem_release_bits_payload_data = {5{$random}};
  assign io_mem_release_bits_payload_client_xact_id = {1{$random}};
  assign io_mem_release_bits_payload_addr = {1{$random}};
//  assign io_mem_release_bits_header_dst = {1{$random}};
//  assign io_mem_release_bits_header_src = {1{$random}};
  assign io_mem_release_valid = 1'h0;
  assign io_mem_probe_ready = 1'h0;
  assign io_mem_finish_bits_payload_manager_xact_id = mem_gxid;
  assign T145 = io_mem_grant_valid ? io_mem_grant_bits_payload_manager_xact_id : mem_gxid;
  assign io_mem_finish_bits_header_dst = mem_gsrc;
  assign T146 = io_mem_grant_valid ? io_mem_grant_bits_header_src : mem_gsrc;
//  assign io_mem_finish_bits_header_src = {1{$random}};
  assign io_mem_finish_valid = T147;
  assign T147 = T151 & mem_needs_ack;
  assign T148 = io_mem_grant_valid ? T149 : mem_needs_ack;
  assign T149 = io_mem_grant_bits_payload_uncached | T150;
  assign T150 = io_mem_grant_bits_payload_g_type != 2'h0;
  assign T151 = state == 4'h7;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_payload_subblock = T152;
  assign T152 = T155 ? T154 : T153;
  assign T153 = 129'hf;
  assign T154 = 129'h3;
  assign T155 = cmd == 4'h1;
  assign io_mem_acquire_bits_payload_a_type = T156;
  assign T156 = T155 ? T158 : T157;
  assign T157 = 2'h0;
  assign T158 = 2'h1;
  assign io_mem_acquire_bits_payload_uncached = T159;
  assign T159 = T155 ? T161 : T160;
  assign T160 = 1'h1;
  assign T161 = 1'h1;
  assign io_mem_acquire_bits_payload_data = T162;
  assign T162 = T163;
  assign T163 = {T168, T164};
  assign T164 = {4'h0, T165};
  assign T165 = mem_req_data[6'h3f:1'h0];
  assign mem_req_data = {T167, T166};
  assign T166 = packet_ram[T137];
  assign T167 = packet_ram[T132];
  assign T168 = {4'h0, T169};
  assign T169 = mem_req_data[7'h7f:7'h40];
  assign io_mem_acquire_bits_payload_client_xact_id = T170;
  assign T170 = T155 ? T172 : T171;
  assign T171 = 2'h0;
  assign T172 = 2'h0;
  assign io_mem_acquire_bits_payload_addr = T173;
  assign T173 = T155 ? T176 : T174;
  assign T174 = T348;
  assign T348 = init_addr[5'h19:1'h0];
  assign init_addr = T175 >> 2'h3;
  assign T175 = addr;
  assign T176 = T349;
  assign T349 = init_addr[5'h19:1'h0];
  assign io_mem_acquire_bits_header_dst = 2'h0;
  assign io_mem_acquire_bits_header_src = 2'h2;
  assign io_mem_acquire_valid = T177;
  assign T177 = T179 | T178;
  assign T178 = state == 4'h4;
  assign T179 = state == 4'h3;
//  assign io_cpu_0_ipi_rep_bits = {1{$random}};
  assign io_cpu_0_ipi_rep_valid = R180;
  assign T350 = reset ? 1'h0 : T181;
  assign T181 = T183 ? 1'h1 : T182;
  assign T182 = io_cpu_0_ipi_rep_ready ? 1'h0 : R180;
  assign T183 = io_cpu_0_ipi_req_valid & T184;
  assign T184 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = pcr_wdata;
  assign io_cpu_0_pcr_req_bits_addr = pcr_addr;
  assign io_cpu_0_pcr_req_bits_rw = T185;
  assign T185 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T186;
  assign T186 = T188 & T187;
  assign T187 = pcr_addr != 5'h1d;
  assign T188 = T189 & T127;
  assign T189 = state == 4'h1;
//  assign io_cpu_0_id = {1{$random}};
  assign io_cpu_0_reset = R190;
  assign T351 = reset ? 1'h1 : T191;
  assign T191 = T193 ? T192 : R190;
  assign T192 = pcr_wdata[1'h0:1'h0];
  assign T193 = T124 & T194;
  assign T194 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T352;
  assign T352 = T195[4'hf:1'h0];
  assign T195 = tx_data >> T196;
  assign T196 = {T197, 4'h0};
  assign T197 = tx_count[1'h1:1'h0];
  assign tx_data = T337 ? tx_header : T198;
  assign T198 = T330 ? pcrReadData : T199;
  assign T199 = packet_ram[packet_ram_raddr];
  assign T200 = T129 ? T203 : T201;
  assign T201 = io_cpu_0_pcr_rep_valid ? io_cpu_0_pcr_rep_bits : T202;
  assign T202 = T124 ? T353 : pcrReadData;
  assign T353 = {63'h0, R190};
  assign T203 = T329 ? T267 : T204;
  assign T204 = T266 ? T236 : T205;
  assign T205 = T235 ? T221 : T206;
  assign T206 = T220 ? T214 : T207;
  assign T207 = T213 ? T211 : T208;
  assign T208 = T209 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T209 = T210[1'h0:1'h0];
  assign T210 = scr_addr;
  assign T211 = T212 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T212 = T210[1'h0:1'h0];
  assign T213 = T210[1'h1:1'h1];
  assign T214 = T219 ? T217 : T215;
  assign T215 = T216 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T216 = T210[1'h0:1'h0];
  assign T217 = T218 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T218 = T210[1'h0:1'h0];
  assign T219 = T210[1'h1:1'h1];
  assign T220 = T210[2'h2:2'h2];
  assign T221 = T234 ? T228 : T222;
  assign T222 = T227 ? T225 : T223;
  assign T223 = T224 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T224 = T210[1'h0:1'h0];
  assign T225 = T226 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T226 = T210[1'h0:1'h0];
  assign T227 = T210[1'h1:1'h1];
  assign T228 = T233 ? T231 : T229;
  assign T229 = T230 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T230 = T210[1'h0:1'h0];
  assign T231 = T232 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T232 = T210[1'h0:1'h0];
  assign T233 = T210[1'h1:1'h1];
  assign T234 = T210[2'h2:2'h2];
  assign T235 = T210[2'h3:2'h3];
  assign T236 = T265 ? T251 : T237;
  assign T237 = T250 ? T244 : T238;
  assign T238 = T243 ? T241 : T239;
  assign T239 = T240 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T240 = T210[1'h0:1'h0];
  assign T241 = T242 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T242 = T210[1'h0:1'h0];
  assign T243 = T210[1'h1:1'h1];
  assign T244 = T249 ? T247 : T245;
  assign T245 = T246 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T246 = T210[1'h0:1'h0];
  assign T247 = T248 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T248 = T210[1'h0:1'h0];
  assign T249 = T210[1'h1:1'h1];
  assign T250 = T210[2'h2:2'h2];
  assign T251 = T264 ? T258 : T252;
  assign T252 = T257 ? T255 : T253;
  assign T253 = T254 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T254 = T210[1'h0:1'h0];
  assign T255 = T256 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T256 = T210[1'h0:1'h0];
  assign T257 = T210[1'h1:1'h1];
  assign T258 = T263 ? T261 : T259;
  assign T259 = T260 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T260 = T210[1'h0:1'h0];
  assign T261 = T262 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T262 = T210[1'h0:1'h0];
  assign T263 = T210[1'h1:1'h1];
  assign T264 = T210[2'h2:2'h2];
  assign T265 = T210[2'h3:2'h3];
  assign T266 = T210[3'h4:3'h4];
  assign T267 = T328 ? T298 : T268;
  assign T268 = T297 ? T283 : T269;
  assign T269 = T282 ? T276 : T270;
  assign T270 = T275 ? T273 : T271;
  assign T271 = T272 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T272 = T210[1'h0:1'h0];
  assign T273 = T274 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T274 = T210[1'h0:1'h0];
  assign T275 = T210[1'h1:1'h1];
  assign T276 = T281 ? T279 : T277;
  assign T277 = T278 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T278 = T210[1'h0:1'h0];
  assign T279 = T280 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T280 = T210[1'h0:1'h0];
  assign T281 = T210[1'h1:1'h1];
  assign T282 = T210[2'h2:2'h2];
  assign T283 = T296 ? T290 : T284;
  assign T284 = T289 ? T287 : T285;
  assign T285 = T286 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T286 = T210[1'h0:1'h0];
  assign T287 = T288 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T288 = T210[1'h0:1'h0];
  assign T289 = T210[1'h1:1'h1];
  assign T290 = T295 ? T293 : T291;
  assign T291 = T292 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T292 = T210[1'h0:1'h0];
  assign T293 = T294 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T294 = T210[1'h0:1'h0];
  assign T295 = T210[1'h1:1'h1];
  assign T296 = T210[2'h2:2'h2];
  assign T297 = T210[2'h3:2'h3];
  assign T298 = T327 ? T313 : T299;
  assign T299 = T312 ? T306 : T300;
  assign T300 = T305 ? T303 : T301;
  assign T301 = T302 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T302 = T210[1'h0:1'h0];
  assign T303 = T304 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T304 = T210[1'h0:1'h0];
  assign T305 = T210[1'h1:1'h1];
  assign T306 = T311 ? T309 : T307;
  assign T307 = T308 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T308 = T210[1'h0:1'h0];
  assign T309 = T310 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T310 = T210[1'h0:1'h0];
  assign T311 = T210[1'h1:1'h1];
  assign T312 = T210[2'h2:2'h2];
  assign T313 = T326 ? T320 : T314;
  assign T314 = T319 ? T317 : T315;
  assign T315 = T316 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T316 = T210[1'h0:1'h0];
  assign T317 = T318 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T318 = T210[1'h0:1'h0];
  assign T319 = T210[1'h1:1'h1];
  assign T320 = T325 ? T323 : T321;
  assign T321 = T322 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T322 = T210[1'h0:1'h0];
  assign T323 = T324 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T324 = T210[1'h0:1'h0];
  assign T325 = T210[1'h1:1'h1];
  assign T326 = T210[2'h2:2'h2];
  assign T327 = T210[2'h3:2'h3];
  assign T328 = T210[3'h4:3'h4];
  assign T329 = T210[3'h5:3'h5];
  assign T330 = T332 | T331;
  assign T331 = cmd == 4'h3;
  assign T332 = cmd == 4'h2;
  assign tx_header = {T334, T333};
  assign T333 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T334 = {addr, seqno};
  assign T335 = T24 ? T336 : seqno;
  assign T336 = rx_shifter_in[5'h17:5'h10];
  assign T337 = tx_word_count == 13'h0;
  assign io_host_out_valid = T338;
  assign T338 = state == 4'h8;
  assign io_host_in_ready = T339;
  assign T339 = state == 4'h0;
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};

  always @(posedge clk) begin
    if (T5)
      packet_ram[T132] <= T1;
    if(reset) begin
      state <= 4'h0;
    end else if(T129) begin
      state <= 4'h8;
    end else if(io_cpu_0_pcr_rep_valid) begin
      state <= 4'h8;
    end else if(T124) begin
      state <= 4'h8;
    end else if(T123) begin
      state <= 4'h2;
    end else if(T113) begin
      state <= T109;
    end else if(T107) begin
      state <= T99;
    end else if(T97) begin
      state <= 4'h7;
    end else if(T92) begin
      state <= 4'h7;
    end else if(T90) begin
      state <= 4'h5;
    end else if(T80) begin
      state <= 4'h6;
    end else if(T67) begin
      state <= T18;
    end
    if(T24) begin
      cmd <= next_cmd;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T29) begin
      rx_count <= 15'h0;
    end else if(T62) begin
      rx_count <= T28;
    end
    if(T24) begin
      size <= T32;
    end
    if(T62) begin
      rx_shifter <= rx_shifter_in;
    end
    if(T107) begin
      addr <= T52;
    end else if(T24) begin
      addr <= T51;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T29) begin
      tx_count <= 15'h0;
    end else if(T61) begin
      tx_count <= T60;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T84) begin
      cnt <= T83;
    end
    if(reset) begin
      mem_acked <= 1'h0;
    end else if(T97) begin
      mem_acked <= 1'h0;
    end else if(T92) begin
      mem_acked <= 1'h0;
    end else if(io_mem_grant_valid) begin
      mem_acked <= 1'h1;
    end
    if(T107) begin
      pos <= T105;
    end else if(T24) begin
      pos <= T104;
    end
    if (T135)
      packet_ram[T137] <= T134;
    if (T139)
      packet_ram[T140] <= rx_shifter_in;
    if(io_mem_grant_valid) begin
      mem_gxid <= io_mem_grant_bits_payload_manager_xact_id;
    end
    if(io_mem_grant_valid) begin
      mem_gsrc <= io_mem_grant_bits_header_src;
    end
    if(io_mem_grant_valid) begin
      mem_needs_ack <= T149;
    end
    if(reset) begin
      R180 <= 1'h0;
    end else if(T183) begin
      R180 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R180 <= 1'h0;
    end
    if(reset) begin
      R190 <= 1'h1;
    end else if(T193) begin
      R190 <= T192;
    end
    if(T129) begin
      pcrReadData <= T203;
    end else if(io_cpu_0_pcr_rep_valid) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T124) begin
      pcrReadData <= T353;
    end
    if(T24) begin
      seqno <= T336;
    end
  end
endmodule

module LockingRRArbiter_9(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [135:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [128:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [135:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [128:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [135:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [128:0] io_in_0_bits_payload_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[135:0] io_out_bits_payload_data,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_a_type,
    output[128:0] io_out_bits_payload_subblock,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T105;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T106;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  reg  locked;
  wire T107;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  reg [1:0] R28;
  wire[1:0] T108;
  wire[1:0] T29;
  wire[128:0] T30;
  wire[128:0] T31;
  wire T32;
  wire[1:0] T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[135:0] T43;
  wire[135:0] T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[25:0] T51;
  wire[25:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire T57;
  wire T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R28 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T105 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T106 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T22 & T18;
  assign T18 = io_out_bits_payload_uncached ? T19 : 1'h0;
  assign T19 = T21 | T20;
  assign T20 = 2'h2 == io_out_bits_payload_a_type;
  assign T21 = 2'h1 == io_out_bits_payload_a_type;
  assign T22 = io_out_ready & io_out_valid;
  assign T107 = reset ? 1'h0 : T23;
  assign T23 = T25 ? 1'h0 : T24;
  assign T24 = T15 ? 1'h1 : locked;
  assign T25 = T22 & T26;
  assign T26 = T27 == 2'h0;
  assign T27 = R28 + 2'h1;
  assign T108 = reset ? 2'h0 : T29;
  assign T29 = T17 ? T27 : R28;
  assign io_out_bits_payload_subblock = T30;
  assign T30 = T34 ? io_in_2_bits_payload_subblock : T31;
  assign T31 = T32 ? io_in_1_bits_payload_subblock : io_in_0_bits_payload_subblock;
  assign T32 = T33[1'h0:1'h0];
  assign T33 = chosen;
  assign T34 = T33[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T35;
  assign T35 = T38 ? io_in_2_bits_payload_a_type : T36;
  assign T36 = T37 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T37 = T33[1'h0:1'h0];
  assign T38 = T33[1'h1:1'h1];
  assign io_out_bits_payload_uncached = T39;
  assign T39 = T42 ? io_in_2_bits_payload_uncached : T40;
  assign T40 = T41 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T41 = T33[1'h0:1'h0];
  assign T42 = T33[1'h1:1'h1];
  assign io_out_bits_payload_data = T43;
  assign T43 = T46 ? io_in_2_bits_payload_data : T44;
  assign T44 = T45 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T45 = T33[1'h0:1'h0];
  assign T46 = T33[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T47;
  assign T47 = T50 ? io_in_2_bits_payload_client_xact_id : T48;
  assign T48 = T49 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T49 = T33[1'h0:1'h0];
  assign T50 = T33[1'h1:1'h1];
  assign io_out_bits_payload_addr = T51;
  assign T51 = T54 ? io_in_2_bits_payload_addr : T52;
  assign T52 = T53 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T53 = T33[1'h0:1'h0];
  assign T54 = T33[1'h1:1'h1];
  assign io_out_bits_header_dst = T55;
  assign T55 = T58 ? io_in_2_bits_header_dst : T56;
  assign T56 = T57 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T57 = T33[1'h0:1'h0];
  assign T58 = T33[1'h1:1'h1];
  assign io_out_bits_header_src = T59;
  assign T59 = T62 ? io_in_2_bits_header_src : T60;
  assign T60 = T61 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T61 = T33[1'h0:1'h0];
  assign T62 = T33[1'h1:1'h1];
  assign io_out_valid = T63;
  assign T63 = T66 ? io_in_2_valid : T64;
  assign T64 = T65 ? io_in_1_valid : io_in_0_valid;
  assign T65 = T33[1'h0:1'h0];
  assign T66 = T33[1'h1:1'h1];
  assign io_in_0_ready = T67;
  assign T67 = T68 & io_out_ready;
  assign T68 = locked ? T80 : T69;
  assign T69 = T79 | T70;
  assign T70 = T71 ^ 1'h1;
  assign T71 = T74 | T72;
  assign T72 = io_in_2_valid & T73;
  assign T73 = last_grant < 2'h2;
  assign T74 = T77 | T75;
  assign T75 = io_in_1_valid & T76;
  assign T76 = last_grant < 2'h1;
  assign T77 = io_in_0_valid & T78;
  assign T78 = last_grant < 2'h0;
  assign T79 = last_grant < 2'h0;
  assign T80 = lockIdx == 2'h0;
  assign io_in_1_ready = T81;
  assign T81 = T82 & io_out_ready;
  assign T82 = locked ? T91 : T83;
  assign T83 = T88 | T84;
  assign T84 = T85 ^ 1'h1;
  assign T85 = T86 | io_in_0_valid;
  assign T86 = T87 | T72;
  assign T87 = T77 | T75;
  assign T88 = T90 & T89;
  assign T89 = last_grant < 2'h1;
  assign T90 = T77 ^ 1'h1;
  assign T91 = lockIdx == 2'h1;
  assign io_in_2_ready = T92;
  assign T92 = T93 & io_out_ready;
  assign T93 = locked ? T104 : T94;
  assign T94 = T100 | T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T97 | io_in_1_valid;
  assign T97 = T98 | io_in_0_valid;
  assign T98 = T99 | T72;
  assign T99 = T77 | T75;
  assign T100 = T102 & T101;
  assign T101 = last_grant < 2'h2;
  assign T102 = T103 ^ 1'h1;
  assign T103 = T77 | T75;
  assign T104 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T25) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R28 <= 2'h0;
    end else if(T17) begin
      R28 <= T27;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [135:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [128:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [135:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [128:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [135:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [128:0] io_in_0_bits_payload_subblock,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[135:0] io_out_2_bits_payload_data,
    output io_out_2_bits_payload_uncached,
    output[1:0] io_out_2_bits_payload_a_type,
    output[128:0] io_out_2_bits_payload_subblock,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[135:0] io_out_1_bits_payload_data,
    output io_out_1_bits_payload_uncached,
    output[1:0] io_out_1_bits_payload_a_type,
    output[128:0] io_out_1_bits_payload_subblock,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[135:0] io_out_0_bits_payload_data,
    output io_out_0_bits_payload_uncached,
    output[1:0] io_out_0_bits_payload_a_type,
    output[128:0] io_out_0_bits_payload_subblock
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_9_io_in_2_ready;
  wire LockingRRArbiter_9_io_in_1_ready;
  wire LockingRRArbiter_9_io_in_0_ready;
  wire LockingRRArbiter_9_io_out_valid;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_9_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_9_io_out_bits_payload_data;
  wire LockingRRArbiter_9_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_9_io_out_bits_payload_a_type;
  wire[128:0] LockingRRArbiter_9_io_out_bits_payload_subblock;
  wire LockingRRArbiter_10_io_in_2_ready;
  wire LockingRRArbiter_10_io_in_1_ready;
  wire LockingRRArbiter_10_io_in_0_ready;
  wire LockingRRArbiter_10_io_out_valid;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_10_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_10_io_out_bits_payload_data;
  wire LockingRRArbiter_10_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_10_io_out_bits_payload_a_type;
  wire[128:0] LockingRRArbiter_10_io_out_bits_payload_subblock;
  wire LockingRRArbiter_11_io_in_2_ready;
  wire LockingRRArbiter_11_io_in_1_ready;
  wire LockingRRArbiter_11_io_in_0_ready;
  wire LockingRRArbiter_11_io_out_valid;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_11_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_11_io_out_bits_payload_data;
  wire LockingRRArbiter_11_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_11_io_out_bits_payload_a_type;
  wire[128:0] LockingRRArbiter_11_io_out_bits_payload_subblock;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_subblock = LockingRRArbiter_9_io_out_bits_payload_subblock;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_9_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_uncached = LockingRRArbiter_9_io_out_bits_payload_uncached;
  assign io_out_0_bits_payload_data = LockingRRArbiter_9_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_9_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_9_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_9_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_9_io_out_valid;
  assign io_out_1_bits_payload_subblock = LockingRRArbiter_10_io_out_bits_payload_subblock;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_10_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_uncached = LockingRRArbiter_10_io_out_bits_payload_uncached;
  assign io_out_1_bits_payload_data = LockingRRArbiter_10_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_10_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_10_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_10_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_10_io_out_valid;
  assign io_out_2_bits_payload_subblock = LockingRRArbiter_11_io_out_bits_payload_subblock;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_11_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_uncached = LockingRRArbiter_11_io_out_bits_payload_uncached;
  assign io_out_2_bits_payload_data = LockingRRArbiter_11_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_11_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_11_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_11_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_11_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_11_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_10_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_9_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_11_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_10_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_9_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_11_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_10_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_9_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_9 LockingRRArbiter_9(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_9_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_9_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_9_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_bits_payload_subblock ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_9_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_9_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_9_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_9_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_9_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_9_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_9_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_9_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_9_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  LockingRRArbiter_9 LockingRRArbiter_10(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_10_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_10_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_10_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_bits_payload_subblock ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_10_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_10_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_10_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_10_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_10_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_10_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_10_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_10_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_10_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  LockingRRArbiter_9 LockingRRArbiter_11(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_11_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_11_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_11_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_bits_payload_subblock ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_11_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_11_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_11_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_11_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_11_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_11_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_11_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_11_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_11_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_10(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [135:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [135:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [135:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[135:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T100;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T101;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  reg  locked;
  wire T102;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  reg [1:0] R31;
  wire[1:0] T103;
  wire[1:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire[135:0] T38;
  wire[135:0] T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire[25:0] T46;
  wire[25:0] T47;
  wire T48;
  wire T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R31 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T100 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T101 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T25 & T18;
  assign T18 = T20 | T19;
  assign T19 = 3'h3 == io_out_bits_payload_r_type;
  assign T20 = T22 | T21;
  assign T21 = 3'h2 == io_out_bits_payload_r_type;
  assign T22 = T24 | T23;
  assign T23 = 3'h1 == io_out_bits_payload_r_type;
  assign T24 = 3'h0 == io_out_bits_payload_r_type;
  assign T25 = io_out_ready & io_out_valid;
  assign T102 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h0 : T27;
  assign T27 = T15 ? 1'h1 : locked;
  assign T28 = T25 & T29;
  assign T29 = T30 == 2'h0;
  assign T30 = R31 + 2'h1;
  assign T103 = reset ? 2'h0 : T32;
  assign T32 = T17 ? T30 : R31;
  assign io_out_bits_payload_r_type = T33;
  assign T33 = T37 ? io_in_2_bits_payload_r_type : T34;
  assign T34 = T35 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = chosen;
  assign T37 = T36[1'h1:1'h1];
  assign io_out_bits_payload_data = T38;
  assign T38 = T41 ? io_in_2_bits_payload_data : T39;
  assign T39 = T40 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T40 = T36[1'h0:1'h0];
  assign T41 = T36[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T42;
  assign T42 = T45 ? io_in_2_bits_payload_client_xact_id : T43;
  assign T43 = T44 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign io_out_bits_payload_addr = T46;
  assign T46 = T49 ? io_in_2_bits_payload_addr : T47;
  assign T47 = T48 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T48 = T36[1'h0:1'h0];
  assign T49 = T36[1'h1:1'h1];
  assign io_out_bits_header_dst = T50;
  assign T50 = T53 ? io_in_2_bits_header_dst : T51;
  assign T51 = T52 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign io_out_bits_header_src = T54;
  assign T54 = T57 ? io_in_2_bits_header_src : T55;
  assign T55 = T56 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T36[1'h1:1'h1];
  assign io_out_valid = T58;
  assign T58 = T61 ? io_in_2_valid : T59;
  assign T59 = T60 ? io_in_1_valid : io_in_0_valid;
  assign T60 = T36[1'h0:1'h0];
  assign T61 = T36[1'h1:1'h1];
  assign io_in_0_ready = T62;
  assign T62 = T63 & io_out_ready;
  assign T63 = locked ? T75 : T64;
  assign T64 = T74 | T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T69 | T67;
  assign T67 = io_in_2_valid & T68;
  assign T68 = last_grant < 2'h2;
  assign T69 = T72 | T70;
  assign T70 = io_in_1_valid & T71;
  assign T71 = last_grant < 2'h1;
  assign T72 = io_in_0_valid & T73;
  assign T73 = last_grant < 2'h0;
  assign T74 = last_grant < 2'h0;
  assign T75 = lockIdx == 2'h0;
  assign io_in_1_ready = T76;
  assign T76 = T77 & io_out_ready;
  assign T77 = locked ? T86 : T78;
  assign T78 = T83 | T79;
  assign T79 = T80 ^ 1'h1;
  assign T80 = T81 | io_in_0_valid;
  assign T81 = T82 | T67;
  assign T82 = T72 | T70;
  assign T83 = T85 & T84;
  assign T84 = last_grant < 2'h1;
  assign T85 = T72 ^ 1'h1;
  assign T86 = lockIdx == 2'h1;
  assign io_in_2_ready = T87;
  assign T87 = T88 & io_out_ready;
  assign T88 = locked ? T99 : T89;
  assign T89 = T95 | T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = T92 | io_in_1_valid;
  assign T92 = T93 | io_in_0_valid;
  assign T93 = T94 | T67;
  assign T94 = T72 | T70;
  assign T95 = T97 & T96;
  assign T96 = last_grant < 2'h2;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T72 | T70;
  assign T99 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T28) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R31 <= 2'h0;
    end else if(T17) begin
      R31 <= T30;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [135:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [135:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [135:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[135:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_r_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[135:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_r_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[135:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_r_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_12_io_in_2_ready;
  wire LockingRRArbiter_12_io_in_1_ready;
  wire LockingRRArbiter_12_io_in_0_ready;
  wire LockingRRArbiter_12_io_out_valid;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_12_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_12_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_12_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_12_io_out_bits_payload_r_type;
  wire LockingRRArbiter_13_io_in_2_ready;
  wire LockingRRArbiter_13_io_in_1_ready;
  wire LockingRRArbiter_13_io_in_0_ready;
  wire LockingRRArbiter_13_io_out_valid;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_13_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_13_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_13_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_13_io_out_bits_payload_r_type;
  wire LockingRRArbiter_14_io_in_2_ready;
  wire LockingRRArbiter_14_io_in_1_ready;
  wire LockingRRArbiter_14_io_in_0_ready;
  wire LockingRRArbiter_14_io_out_valid;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_14_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_14_io_out_bits_payload_client_xact_id;
  wire[135:0] LockingRRArbiter_14_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_14_io_out_bits_payload_r_type;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_12_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_12_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_12_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_12_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_12_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_12_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_12_io_out_valid;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_13_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_13_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_13_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_13_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_13_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_13_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_13_io_out_valid;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_14_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_14_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_14_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_14_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_14_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_14_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_14_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_14_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_13_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_12_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_14_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_13_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_12_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_14_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_13_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_12_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_10 LockingRRArbiter_12(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_12_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_12_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_12_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_12_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_12_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_12_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_12_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_12_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_12_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_12_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_10 LockingRRArbiter_13(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_13_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_13_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_13_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_13_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_13_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_13_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_13_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_13_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_13_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_13_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_10 LockingRRArbiter_14(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_14_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_14_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_14_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_14_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_14_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_14_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_14_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_14_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_14_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_14_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_11(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_p_type,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T62;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[25:0] T14;
  wire[25:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T62 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_payload_p_type = T9;
  assign T9 = T13 ? io_in_2_bits_payload_p_type : T10;
  assign T10 = T11 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1:1'h1];
  assign io_out_bits_payload_addr = T14;
  assign T14 = T17 ? io_in_2_bits_payload_addr : T15;
  assign T15 = T16 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T16 = T12[1'h0:1'h0];
  assign T17 = T12[1'h1:1'h1];
  assign io_out_bits_header_dst = T18;
  assign T18 = T21 ? io_in_2_bits_header_dst : T19;
  assign T19 = T20 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign io_out_bits_header_src = T22;
  assign T22 = T25 ? io_in_2_bits_header_src : T23;
  assign T23 = T24 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T12[1'h1:1'h1];
  assign io_out_valid = T26;
  assign T26 = T29 ? io_in_2_valid : T27;
  assign T27 = T28 ? io_in_1_valid : io_in_0_valid;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign io_in_0_ready = T30;
  assign T30 = T31 & io_out_ready;
  assign T31 = T41 | T32;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T36 | T34;
  assign T34 = io_in_2_valid & T35;
  assign T35 = last_grant < 2'h2;
  assign T36 = T39 | T37;
  assign T37 = io_in_1_valid & T38;
  assign T38 = last_grant < 2'h1;
  assign T39 = io_in_0_valid & T40;
  assign T40 = last_grant < 2'h0;
  assign T41 = last_grant < 2'h0;
  assign io_in_1_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = T48 | T44;
  assign T44 = T45 ^ 1'h1;
  assign T45 = T46 | io_in_0_valid;
  assign T46 = T47 | T34;
  assign T47 = T39 | T37;
  assign T48 = T50 & T49;
  assign T49 = last_grant < 2'h1;
  assign T50 = T39 ^ 1'h1;
  assign io_in_2_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T58 | T53;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T55 | io_in_1_valid;
  assign T55 = T56 | io_in_0_valid;
  assign T56 = T57 | T34;
  assign T57 = T39 | T37;
  assign T58 = T60 & T59;
  assign T59 = last_grant < 2'h2;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T39 | T37;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_15_io_in_2_ready;
  wire LockingRRArbiter_15_io_in_1_ready;
  wire LockingRRArbiter_15_io_in_0_ready;
  wire LockingRRArbiter_15_io_out_valid;
  wire[1:0] LockingRRArbiter_15_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_15_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_15_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_15_io_out_bits_payload_p_type;
  wire LockingRRArbiter_16_io_in_2_ready;
  wire LockingRRArbiter_16_io_in_1_ready;
  wire LockingRRArbiter_16_io_in_0_ready;
  wire LockingRRArbiter_16_io_out_valid;
  wire[1:0] LockingRRArbiter_16_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_16_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_16_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_16_io_out_bits_payload_p_type;
  wire LockingRRArbiter_17_io_in_2_ready;
  wire LockingRRArbiter_17_io_in_1_ready;
  wire LockingRRArbiter_17_io_in_0_ready;
  wire LockingRRArbiter_17_io_out_valid;
  wire[1:0] LockingRRArbiter_17_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_17_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_17_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_17_io_out_bits_payload_p_type;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_15_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_15_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_15_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_15_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_15_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_16_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_16_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_16_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_16_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_16_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_17_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_17_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_17_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_17_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_17_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_17_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_16_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_15_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_17_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_16_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_15_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_17_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_16_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_15_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_11 LockingRRArbiter_15(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_15_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_15_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_15_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_15_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_15_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_15_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_15_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( LockingRRArbiter_15_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_11 LockingRRArbiter_16(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_16_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_16_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_16_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_16_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_16_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_16_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_16_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( LockingRRArbiter_16_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_11 LockingRRArbiter_17(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_17_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_17_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_17_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_17_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_17_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_17_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_17_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( LockingRRArbiter_17_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_12(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [135:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [135:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [135:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[135:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T104;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T105;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  reg  locked;
  wire T106;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  reg [1:0] R31;
  wire[1:0] T107;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[3:0] T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire[135:0] T50;
  wire[135:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R31 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T104 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T105 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T25 & T18;
  assign T18 = io_out_bits_payload_uncached ? T22 : T19;
  assign T19 = T21 | T20;
  assign T20 = 2'h2 == io_out_bits_payload_g_type;
  assign T21 = 2'h1 == io_out_bits_payload_g_type;
  assign T22 = T24 | T23;
  assign T23 = 2'h2 == io_out_bits_payload_g_type;
  assign T24 = 2'h0 == io_out_bits_payload_g_type;
  assign T25 = io_out_ready & io_out_valid;
  assign T106 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h0 : T27;
  assign T27 = T15 ? 1'h1 : locked;
  assign T28 = T25 & T29;
  assign T29 = T30 == 2'h0;
  assign T30 = R31 + 2'h1;
  assign T107 = reset ? 2'h0 : T32;
  assign T32 = T17 ? T30 : R31;
  assign io_out_bits_payload_g_type = T33;
  assign T33 = T37 ? io_in_2_bits_payload_g_type : T34;
  assign T34 = T35 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = chosen;
  assign T37 = T36[1'h1:1'h1];
  assign io_out_bits_payload_uncached = T38;
  assign T38 = T41 ? io_in_2_bits_payload_uncached : T39;
  assign T39 = T40 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T40 = T36[1'h0:1'h0];
  assign T41 = T36[1'h1:1'h1];
  assign io_out_bits_payload_manager_xact_id = T42;
  assign T42 = T45 ? io_in_2_bits_payload_manager_xact_id : T43;
  assign T43 = T44 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T46;
  assign T46 = T49 ? io_in_2_bits_payload_client_xact_id : T47;
  assign T47 = T48 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T48 = T36[1'h0:1'h0];
  assign T49 = T36[1'h1:1'h1];
  assign io_out_bits_payload_data = T50;
  assign T50 = T53 ? io_in_2_bits_payload_data : T51;
  assign T51 = T52 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign io_out_bits_header_dst = T54;
  assign T54 = T57 ? io_in_2_bits_header_dst : T55;
  assign T55 = T56 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T36[1'h1:1'h1];
  assign io_out_bits_header_src = T58;
  assign T58 = T61 ? io_in_2_bits_header_src : T59;
  assign T59 = T60 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T60 = T36[1'h0:1'h0];
  assign T61 = T36[1'h1:1'h1];
  assign io_out_valid = T62;
  assign T62 = T65 ? io_in_2_valid : T63;
  assign T63 = T64 ? io_in_1_valid : io_in_0_valid;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T36[1'h1:1'h1];
  assign io_in_0_ready = T66;
  assign T66 = T67 & io_out_ready;
  assign T67 = locked ? T79 : T68;
  assign T68 = T78 | T69;
  assign T69 = T70 ^ 1'h1;
  assign T70 = T73 | T71;
  assign T71 = io_in_2_valid & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T76 | T74;
  assign T74 = io_in_1_valid & T75;
  assign T75 = last_grant < 2'h1;
  assign T76 = io_in_0_valid & T77;
  assign T77 = last_grant < 2'h0;
  assign T78 = last_grant < 2'h0;
  assign T79 = lockIdx == 2'h0;
  assign io_in_1_ready = T80;
  assign T80 = T81 & io_out_ready;
  assign T81 = locked ? T90 : T82;
  assign T82 = T87 | T83;
  assign T83 = T84 ^ 1'h1;
  assign T84 = T85 | io_in_0_valid;
  assign T85 = T86 | T71;
  assign T86 = T76 | T74;
  assign T87 = T89 & T88;
  assign T88 = last_grant < 2'h1;
  assign T89 = T76 ^ 1'h1;
  assign T90 = lockIdx == 2'h1;
  assign io_in_2_ready = T91;
  assign T91 = T92 & io_out_ready;
  assign T92 = locked ? T103 : T93;
  assign T93 = T99 | T94;
  assign T94 = T95 ^ 1'h1;
  assign T95 = T96 | io_in_1_valid;
  assign T96 = T97 | io_in_0_valid;
  assign T97 = T98 | T71;
  assign T98 = T76 | T74;
  assign T99 = T101 & T100;
  assign T100 = last_grant < 2'h2;
  assign T101 = T102 ^ 1'h1;
  assign T102 = T76 | T74;
  assign T103 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T28) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R31 <= 2'h0;
    end else if(T17) begin
      R31 <= T30;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [135:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [135:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [135:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[135:0] io_out_2_bits_payload_data,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[3:0] io_out_2_bits_payload_manager_xact_id,
    output io_out_2_bits_payload_uncached,
    output[1:0] io_out_2_bits_payload_g_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[135:0] io_out_1_bits_payload_data,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[3:0] io_out_1_bits_payload_manager_xact_id,
    output io_out_1_bits_payload_uncached,
    output[1:0] io_out_1_bits_payload_g_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[135:0] io_out_0_bits_payload_data,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[3:0] io_out_0_bits_payload_manager_xact_id,
    output io_out_0_bits_payload_uncached,
    output[1:0] io_out_0_bits_payload_g_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_18_io_in_2_ready;
  wire LockingRRArbiter_18_io_in_1_ready;
  wire LockingRRArbiter_18_io_in_0_ready;
  wire LockingRRArbiter_18_io_out_valid;
  wire[1:0] LockingRRArbiter_18_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_18_io_out_bits_header_dst;
  wire[135:0] LockingRRArbiter_18_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_18_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_18_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_18_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_18_io_out_bits_payload_g_type;
  wire LockingRRArbiter_19_io_in_2_ready;
  wire LockingRRArbiter_19_io_in_1_ready;
  wire LockingRRArbiter_19_io_in_0_ready;
  wire LockingRRArbiter_19_io_out_valid;
  wire[1:0] LockingRRArbiter_19_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_19_io_out_bits_header_dst;
  wire[135:0] LockingRRArbiter_19_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_19_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_19_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_19_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_19_io_out_bits_payload_g_type;
  wire LockingRRArbiter_20_io_in_2_ready;
  wire LockingRRArbiter_20_io_in_1_ready;
  wire LockingRRArbiter_20_io_in_0_ready;
  wire LockingRRArbiter_20_io_out_valid;
  wire[1:0] LockingRRArbiter_20_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_20_io_out_bits_header_dst;
  wire[135:0] LockingRRArbiter_20_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_20_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_20_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_20_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_20_io_out_bits_payload_g_type;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_18_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_uncached = LockingRRArbiter_18_io_out_bits_payload_uncached;
  assign io_out_0_bits_payload_manager_xact_id = LockingRRArbiter_18_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_18_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_data = LockingRRArbiter_18_io_out_bits_payload_data;
  assign io_out_0_bits_header_dst = LockingRRArbiter_18_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_18_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_18_io_out_valid;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_19_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_uncached = LockingRRArbiter_19_io_out_bits_payload_uncached;
  assign io_out_1_bits_payload_manager_xact_id = LockingRRArbiter_19_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_19_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_data = LockingRRArbiter_19_io_out_bits_payload_data;
  assign io_out_1_bits_header_dst = LockingRRArbiter_19_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_19_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_19_io_out_valid;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_20_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_uncached = LockingRRArbiter_20_io_out_bits_payload_uncached;
  assign io_out_2_bits_payload_manager_xact_id = LockingRRArbiter_20_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_20_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_data = LockingRRArbiter_20_io_out_bits_payload_data;
  assign io_out_2_bits_header_dst = LockingRRArbiter_20_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_20_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_20_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_20_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_19_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_18_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_20_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_19_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_18_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_20_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_19_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_18_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_12 LockingRRArbiter_18(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_18_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_18_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_18_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_18_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_18_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_18_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_18_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_18_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_18_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_18_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_18_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_12 LockingRRArbiter_19(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_19_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_19_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_19_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_19_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_19_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_19_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_19_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_19_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_19_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_19_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_19_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_12 LockingRRArbiter_20(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_20_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_uncached( io_in_2_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_20_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_uncached( io_in_1_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_20_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_uncached( io_in_0_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_20_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_20_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_20_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_20_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_20_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_20_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_20_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_20_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_13(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T58;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T58 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_payload_manager_xact_id = T9;
  assign T9 = T13 ? io_in_2_bits_payload_manager_xact_id : T10;
  assign T10 = T11 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1:1'h1];
  assign io_out_bits_header_dst = T14;
  assign T14 = T17 ? io_in_2_bits_header_dst : T15;
  assign T15 = T16 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T16 = T12[1'h0:1'h0];
  assign T17 = T12[1'h1:1'h1];
  assign io_out_bits_header_src = T18;
  assign T18 = T21 ? io_in_2_bits_header_src : T19;
  assign T19 = T20 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign io_out_valid = T22;
  assign T22 = T25 ? io_in_2_valid : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T12[1'h1:1'h1];
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T37 | T28;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T32 | T30;
  assign T30 = io_in_2_valid & T31;
  assign T31 = last_grant < 2'h2;
  assign T32 = T35 | T33;
  assign T33 = io_in_1_valid & T34;
  assign T34 = last_grant < 2'h1;
  assign T35 = io_in_0_valid & T36;
  assign T36 = last_grant < 2'h0;
  assign T37 = last_grant < 2'h0;
  assign io_in_1_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T44 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T42 | io_in_0_valid;
  assign T42 = T43 | T30;
  assign T43 = T35 | T33;
  assign T44 = T46 & T45;
  assign T45 = last_grant < 2'h1;
  assign T46 = T35 ^ 1'h1;
  assign io_in_2_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T54 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_1_valid;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T30;
  assign T53 = T35 | T33;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h2;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T35 | T33;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[3:0] io_out_2_bits_payload_manager_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[3:0] io_out_1_bits_payload_manager_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[3:0] io_out_0_bits_payload_manager_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_21_io_in_2_ready;
  wire LockingRRArbiter_21_io_in_1_ready;
  wire LockingRRArbiter_21_io_in_0_ready;
  wire LockingRRArbiter_21_io_out_valid;
  wire[1:0] LockingRRArbiter_21_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_21_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_21_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_22_io_in_2_ready;
  wire LockingRRArbiter_22_io_in_1_ready;
  wire LockingRRArbiter_22_io_in_0_ready;
  wire LockingRRArbiter_22_io_out_valid;
  wire[1:0] LockingRRArbiter_22_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_22_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_22_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_23_io_in_2_ready;
  wire LockingRRArbiter_23_io_in_1_ready;
  wire LockingRRArbiter_23_io_in_0_ready;
  wire LockingRRArbiter_23_io_out_valid;
  wire[1:0] LockingRRArbiter_23_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_23_io_out_bits_header_dst;
  wire[3:0] LockingRRArbiter_23_io_out_bits_payload_manager_xact_id;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_manager_xact_id = LockingRRArbiter_21_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_21_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_21_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_21_io_out_valid;
  assign io_out_1_bits_payload_manager_xact_id = LockingRRArbiter_22_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_22_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_22_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_22_io_out_valid;
  assign io_out_2_bits_payload_manager_xact_id = LockingRRArbiter_23_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_23_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_23_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_23_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_23_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_22_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_21_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_23_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_22_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_21_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_23_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_22_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_21_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_13 LockingRRArbiter_21(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_21_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_21_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_21_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_21_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_21_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_21_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_21_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_13 LockingRRArbiter_22(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_22_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_22_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_22_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_22_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_22_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_22_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_22_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_13 LockingRRArbiter_23(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_23_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_bits_payload_manager_xact_id ),
       .io_in_1_ready( LockingRRArbiter_23_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_bits_payload_manager_xact_id ),
       .io_in_0_ready( LockingRRArbiter_23_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_23_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_23_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_23_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_23_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketChipCrossbarNetwork(input clk, input reset,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [1:0] io_clients_1_acquire_bits_header_src,
    input [1:0] io_clients_1_acquire_bits_header_dst,
    input [25:0] io_clients_1_acquire_bits_payload_addr,
    input [1:0] io_clients_1_acquire_bits_payload_client_xact_id,
    input [135:0] io_clients_1_acquire_bits_payload_data,
    input  io_clients_1_acquire_bits_payload_uncached,
    input [1:0] io_clients_1_acquire_bits_payload_a_type,
    input [128:0] io_clients_1_acquire_bits_payload_subblock,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_header_src,
    output[1:0] io_clients_1_grant_bits_header_dst,
    output[135:0] io_clients_1_grant_bits_payload_data,
    output[1:0] io_clients_1_grant_bits_payload_client_xact_id,
    output[3:0] io_clients_1_grant_bits_payload_manager_xact_id,
    output io_clients_1_grant_bits_payload_uncached,
    output[1:0] io_clients_1_grant_bits_payload_g_type,
    output io_clients_1_finish_ready,
    input  io_clients_1_finish_valid,
    input [1:0] io_clients_1_finish_bits_header_src,
    input [1:0] io_clients_1_finish_bits_header_dst,
    input [3:0] io_clients_1_finish_bits_payload_manager_xact_id,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[1:0] io_clients_1_probe_bits_header_src,
    output[1:0] io_clients_1_probe_bits_header_dst,
    output[25:0] io_clients_1_probe_bits_payload_addr,
    output[1:0] io_clients_1_probe_bits_payload_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_header_src,
    input [1:0] io_clients_1_release_bits_header_dst,
    input [25:0] io_clients_1_release_bits_payload_addr,
    input [1:0] io_clients_1_release_bits_payload_client_xact_id,
    input [135:0] io_clients_1_release_bits_payload_data,
    input [2:0] io_clients_1_release_bits_payload_r_type,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [1:0] io_clients_0_acquire_bits_header_src,
    input [1:0] io_clients_0_acquire_bits_header_dst,
    input [25:0] io_clients_0_acquire_bits_payload_addr,
    input [1:0] io_clients_0_acquire_bits_payload_client_xact_id,
    input [135:0] io_clients_0_acquire_bits_payload_data,
    input  io_clients_0_acquire_bits_payload_uncached,
    input [1:0] io_clients_0_acquire_bits_payload_a_type,
    input [128:0] io_clients_0_acquire_bits_payload_subblock,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_header_src,
    output[1:0] io_clients_0_grant_bits_header_dst,
    output[135:0] io_clients_0_grant_bits_payload_data,
    output[1:0] io_clients_0_grant_bits_payload_client_xact_id,
    output[3:0] io_clients_0_grant_bits_payload_manager_xact_id,
    output io_clients_0_grant_bits_payload_uncached,
    output[1:0] io_clients_0_grant_bits_payload_g_type,
    output io_clients_0_finish_ready,
    input  io_clients_0_finish_valid,
    input [1:0] io_clients_0_finish_bits_header_src,
    input [1:0] io_clients_0_finish_bits_header_dst,
    input [3:0] io_clients_0_finish_bits_payload_manager_xact_id,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[1:0] io_clients_0_probe_bits_header_src,
    output[1:0] io_clients_0_probe_bits_header_dst,
    output[25:0] io_clients_0_probe_bits_payload_addr,
    output[1:0] io_clients_0_probe_bits_payload_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_header_src,
    input [1:0] io_clients_0_release_bits_header_dst,
    input [25:0] io_clients_0_release_bits_payload_addr,
    input [1:0] io_clients_0_release_bits_payload_client_xact_id,
    input [135:0] io_clients_0_release_bits_payload_data,
    input [2:0] io_clients_0_release_bits_payload_r_type,
    input  io_managers_0_acquire_ready,
    output io_managers_0_acquire_valid,
    output[1:0] io_managers_0_acquire_bits_header_src,
    output[1:0] io_managers_0_acquire_bits_header_dst,
    output[25:0] io_managers_0_acquire_bits_payload_addr,
    output[1:0] io_managers_0_acquire_bits_payload_client_xact_id,
    output[135:0] io_managers_0_acquire_bits_payload_data,
    output io_managers_0_acquire_bits_payload_uncached,
    output[1:0] io_managers_0_acquire_bits_payload_a_type,
    output[128:0] io_managers_0_acquire_bits_payload_subblock,
    output io_managers_0_grant_ready,
    input  io_managers_0_grant_valid,
    input [1:0] io_managers_0_grant_bits_header_src,
    input [1:0] io_managers_0_grant_bits_header_dst,
    input [135:0] io_managers_0_grant_bits_payload_data,
    input [1:0] io_managers_0_grant_bits_payload_client_xact_id,
    input [3:0] io_managers_0_grant_bits_payload_manager_xact_id,
    input  io_managers_0_grant_bits_payload_uncached,
    input [1:0] io_managers_0_grant_bits_payload_g_type,
    input  io_managers_0_finish_ready,
    output io_managers_0_finish_valid,
    output[1:0] io_managers_0_finish_bits_header_src,
    output[1:0] io_managers_0_finish_bits_header_dst,
    output[3:0] io_managers_0_finish_bits_payload_manager_xact_id,
    output io_managers_0_probe_ready,
    input  io_managers_0_probe_valid,
    input [1:0] io_managers_0_probe_bits_header_src,
    input [1:0] io_managers_0_probe_bits_header_dst,
    input [25:0] io_managers_0_probe_bits_payload_addr,
    input [1:0] io_managers_0_probe_bits_payload_p_type,
    input  io_managers_0_release_ready,
    output io_managers_0_release_valid,
    output[1:0] io_managers_0_release_bits_header_src,
    output[1:0] io_managers_0_release_bits_header_dst,
    output[25:0] io_managers_0_release_bits_payload_addr,
    output[1:0] io_managers_0_release_bits_payload_client_xact_id,
    output[135:0] io_managers_0_release_bits_payload_data,
    output[2:0] io_managers_0_release_bits_payload_r_type
);

  wire T0;
  wire[3:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire[3:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[3:0] T15;
  wire[1:0] T16;
  wire[135:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire[2:0] T31;
  wire[135:0] T32;
  wire[1:0] T33;
  wire[25:0] T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[2:0] T39;
  wire[135:0] T40;
  wire[1:0] T41;
  wire[25:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire[128:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[135:0] T51;
  wire[1:0] T52;
  wire[25:0] T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire T57;
  wire[128:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[135:0] T61;
  wire[1:0] T62;
  wire[25:0] T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire T67;
  wire[2:0] T68;
  wire[135:0] T69;
  wire[1:0] T70;
  wire[25:0] T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire T75;
  wire T76;
  wire[3:0] T77;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire T81;
  wire T82;
  wire[128:0] T83;
  wire[1:0] T84;
  wire T85;
  wire[135:0] T86;
  wire[1:0] T87;
  wire[25:0] T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire T92;
  wire T93;
  wire[1:0] T94;
  wire[25:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire T99;
  wire T100;
  wire[1:0] T101;
  wire T102;
  wire[3:0] T103;
  wire[1:0] T104;
  wire[135:0] T105;
  wire[1:0] T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire T109;
  wire T110;
  wire T111;
  wire[1:0] T112;
  wire[25:0] T113;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire T120;
  wire[3:0] T121;
  wire[1:0] T122;
  wire[135:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire acqNet_io_in_2_ready;
  wire acqNet_io_in_1_ready;
  wire acqNet_io_out_0_valid;
  wire[1:0] acqNet_io_out_0_bits_header_src;
  wire[1:0] acqNet_io_out_0_bits_header_dst;
  wire[25:0] acqNet_io_out_0_bits_payload_addr;
  wire[1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[135:0] acqNet_io_out_0_bits_payload_data;
  wire acqNet_io_out_0_bits_payload_uncached;
  wire[1:0] acqNet_io_out_0_bits_payload_a_type;
  wire[128:0] acqNet_io_out_0_bits_payload_subblock;
  wire relNet_io_in_2_ready;
  wire relNet_io_in_1_ready;
  wire relNet_io_out_0_valid;
  wire[1:0] relNet_io_out_0_bits_header_src;
  wire[1:0] relNet_io_out_0_bits_header_dst;
  wire[25:0] relNet_io_out_0_bits_payload_addr;
  wire[1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire[135:0] relNet_io_out_0_bits_payload_data;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire prbNet_io_in_0_ready;
  wire prbNet_io_out_2_valid;
  wire[1:0] prbNet_io_out_2_bits_header_src;
  wire[1:0] prbNet_io_out_2_bits_header_dst;
  wire[25:0] prbNet_io_out_2_bits_payload_addr;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire prbNet_io_out_1_valid;
  wire[1:0] prbNet_io_out_1_bits_header_src;
  wire[1:0] prbNet_io_out_1_bits_header_dst;
  wire[25:0] prbNet_io_out_1_bits_payload_addr;
  wire[1:0] prbNet_io_out_1_bits_payload_p_type;
  wire gntNet_io_in_0_ready;
  wire gntNet_io_out_2_valid;
  wire[1:0] gntNet_io_out_2_bits_header_src;
  wire[1:0] gntNet_io_out_2_bits_header_dst;
  wire[135:0] gntNet_io_out_2_bits_payload_data;
  wire[1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[3:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire gntNet_io_out_2_bits_payload_uncached;
  wire[1:0] gntNet_io_out_2_bits_payload_g_type;
  wire gntNet_io_out_1_valid;
  wire[1:0] gntNet_io_out_1_bits_header_src;
  wire[1:0] gntNet_io_out_1_bits_header_dst;
  wire[135:0] gntNet_io_out_1_bits_payload_data;
  wire[1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire[3:0] gntNet_io_out_1_bits_payload_manager_xact_id;
  wire gntNet_io_out_1_bits_payload_uncached;
  wire[1:0] gntNet_io_out_1_bits_payload_g_type;
  wire ackNet_io_in_2_ready;
  wire ackNet_io_in_1_ready;
  wire ackNet_io_out_0_valid;
  wire[1:0] ackNet_io_out_0_bits_header_src;
  wire[1:0] ackNet_io_out_0_bits_header_dst;
  wire[3:0] ackNet_io_out_0_bits_payload_manager_xact_id;


  assign T0 = io_managers_0_finish_ready;
  assign T1 = io_clients_0_finish_bits_payload_manager_xact_id;
  assign T2 = io_clients_0_finish_bits_header_dst;
  assign T3 = T4;
  assign T4 = io_clients_0_finish_bits_header_src + 2'h1;
  assign T5 = io_clients_0_finish_valid;
  assign T6 = io_clients_1_finish_bits_payload_manager_xact_id;
  assign T7 = io_clients_1_finish_bits_header_dst;
  assign T8 = T9;
  assign T9 = io_clients_1_finish_bits_header_src + 2'h1;
  assign T10 = io_clients_1_finish_valid;
  assign T11 = io_clients_0_grant_ready;
  assign T12 = io_clients_1_grant_ready;
  assign T13 = io_managers_0_grant_bits_payload_g_type;
  assign T14 = io_managers_0_grant_bits_payload_uncached;
  assign T15 = io_managers_0_grant_bits_payload_manager_xact_id;
  assign T16 = io_managers_0_grant_bits_payload_client_xact_id;
  assign T17 = io_managers_0_grant_bits_payload_data;
  assign T18 = T19;
  assign T19 = io_managers_0_grant_bits_header_dst + 2'h1;
  assign T20 = io_managers_0_grant_bits_header_src;
  assign T21 = io_managers_0_grant_valid;
  assign T22 = io_clients_0_probe_ready;
  assign T23 = io_clients_1_probe_ready;
  assign T24 = io_managers_0_probe_bits_payload_p_type;
  assign T25 = io_managers_0_probe_bits_payload_addr;
  assign T26 = T27;
  assign T27 = io_managers_0_probe_bits_header_dst + 2'h1;
  assign T28 = io_managers_0_probe_bits_header_src;
  assign T29 = io_managers_0_probe_valid;
  assign T30 = io_managers_0_release_ready;
  assign T31 = io_clients_0_release_bits_payload_r_type;
  assign T32 = io_clients_0_release_bits_payload_data;
  assign T33 = io_clients_0_release_bits_payload_client_xact_id;
  assign T34 = io_clients_0_release_bits_payload_addr;
  assign T35 = io_clients_0_release_bits_header_dst;
  assign T36 = T37;
  assign T37 = io_clients_0_release_bits_header_src + 2'h1;
  assign T38 = io_clients_0_release_valid;
  assign T39 = io_clients_1_release_bits_payload_r_type;
  assign T40 = io_clients_1_release_bits_payload_data;
  assign T41 = io_clients_1_release_bits_payload_client_xact_id;
  assign T42 = io_clients_1_release_bits_payload_addr;
  assign T43 = io_clients_1_release_bits_header_dst;
  assign T44 = T45;
  assign T45 = io_clients_1_release_bits_header_src + 2'h1;
  assign T46 = io_clients_1_release_valid;
  assign T47 = io_managers_0_acquire_ready;
  assign T48 = io_clients_0_acquire_bits_payload_subblock;
  assign T49 = io_clients_0_acquire_bits_payload_a_type;
  assign T50 = io_clients_0_acquire_bits_payload_uncached;
  assign T51 = io_clients_0_acquire_bits_payload_data;
  assign T52 = io_clients_0_acquire_bits_payload_client_xact_id;
  assign T53 = io_clients_0_acquire_bits_payload_addr;
  assign T54 = io_clients_0_acquire_bits_header_dst;
  assign T55 = T56;
  assign T56 = io_clients_0_acquire_bits_header_src + 2'h1;
  assign T57 = io_clients_0_acquire_valid;
  assign T58 = io_clients_1_acquire_bits_payload_subblock;
  assign T59 = io_clients_1_acquire_bits_payload_a_type;
  assign T60 = io_clients_1_acquire_bits_payload_uncached;
  assign T61 = io_clients_1_acquire_bits_payload_data;
  assign T62 = io_clients_1_acquire_bits_payload_client_xact_id;
  assign T63 = io_clients_1_acquire_bits_payload_addr;
  assign T64 = io_clients_1_acquire_bits_header_dst;
  assign T65 = T66;
  assign T66 = io_clients_1_acquire_bits_header_src + 2'h1;
  assign T67 = io_clients_1_acquire_valid;
  assign io_managers_0_release_bits_payload_r_type = T68;
  assign T68 = relNet_io_out_0_bits_payload_r_type;
  assign io_managers_0_release_bits_payload_data = T69;
  assign T69 = relNet_io_out_0_bits_payload_data;
  assign io_managers_0_release_bits_payload_client_xact_id = T70;
  assign T70 = relNet_io_out_0_bits_payload_client_xact_id;
  assign io_managers_0_release_bits_payload_addr = T71;
  assign T71 = relNet_io_out_0_bits_payload_addr;
  assign io_managers_0_release_bits_header_dst = T72;
  assign T72 = relNet_io_out_0_bits_header_dst;
  assign io_managers_0_release_bits_header_src = T73;
  assign T73 = T74;
  assign T74 = relNet_io_out_0_bits_header_src - 2'h1;
  assign io_managers_0_release_valid = T75;
  assign T75 = relNet_io_out_0_valid;
  assign io_managers_0_probe_ready = T76;
  assign T76 = prbNet_io_in_0_ready;
  assign io_managers_0_finish_bits_payload_manager_xact_id = T77;
  assign T77 = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign io_managers_0_finish_bits_header_dst = T78;
  assign T78 = ackNet_io_out_0_bits_header_dst;
  assign io_managers_0_finish_bits_header_src = T79;
  assign T79 = T80;
  assign T80 = ackNet_io_out_0_bits_header_src - 2'h1;
  assign io_managers_0_finish_valid = T81;
  assign T81 = ackNet_io_out_0_valid;
  assign io_managers_0_grant_ready = T82;
  assign T82 = gntNet_io_in_0_ready;
  assign io_managers_0_acquire_bits_payload_subblock = T83;
  assign T83 = acqNet_io_out_0_bits_payload_subblock;
  assign io_managers_0_acquire_bits_payload_a_type = T84;
  assign T84 = acqNet_io_out_0_bits_payload_a_type;
  assign io_managers_0_acquire_bits_payload_uncached = T85;
  assign T85 = acqNet_io_out_0_bits_payload_uncached;
  assign io_managers_0_acquire_bits_payload_data = T86;
  assign T86 = acqNet_io_out_0_bits_payload_data;
  assign io_managers_0_acquire_bits_payload_client_xact_id = T87;
  assign T87 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign io_managers_0_acquire_bits_payload_addr = T88;
  assign T88 = acqNet_io_out_0_bits_payload_addr;
  assign io_managers_0_acquire_bits_header_dst = T89;
  assign T89 = acqNet_io_out_0_bits_header_dst;
  assign io_managers_0_acquire_bits_header_src = T90;
  assign T90 = T91;
  assign T91 = acqNet_io_out_0_bits_header_src - 2'h1;
  assign io_managers_0_acquire_valid = T92;
  assign T92 = acqNet_io_out_0_valid;
  assign io_clients_0_release_ready = T93;
  assign T93 = relNet_io_in_1_ready;
  assign io_clients_0_probe_bits_payload_p_type = T94;
  assign T94 = prbNet_io_out_1_bits_payload_p_type;
  assign io_clients_0_probe_bits_payload_addr = T95;
  assign T95 = prbNet_io_out_1_bits_payload_addr;
  assign io_clients_0_probe_bits_header_dst = T96;
  assign T96 = T97;
  assign T97 = prbNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_probe_bits_header_src = T98;
  assign T98 = prbNet_io_out_1_bits_header_src;
  assign io_clients_0_probe_valid = T99;
  assign T99 = prbNet_io_out_1_valid;
  assign io_clients_0_finish_ready = T100;
  assign T100 = ackNet_io_in_1_ready;
  assign io_clients_0_grant_bits_payload_g_type = T101;
  assign T101 = gntNet_io_out_1_bits_payload_g_type;
  assign io_clients_0_grant_bits_payload_uncached = T102;
  assign T102 = gntNet_io_out_1_bits_payload_uncached;
  assign io_clients_0_grant_bits_payload_manager_xact_id = T103;
  assign T103 = gntNet_io_out_1_bits_payload_manager_xact_id;
  assign io_clients_0_grant_bits_payload_client_xact_id = T104;
  assign T104 = gntNet_io_out_1_bits_payload_client_xact_id;
  assign io_clients_0_grant_bits_payload_data = T105;
  assign T105 = gntNet_io_out_1_bits_payload_data;
  assign io_clients_0_grant_bits_header_dst = T106;
  assign T106 = T107;
  assign T107 = gntNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_grant_bits_header_src = T108;
  assign T108 = gntNet_io_out_1_bits_header_src;
  assign io_clients_0_grant_valid = T109;
  assign T109 = gntNet_io_out_1_valid;
  assign io_clients_0_acquire_ready = T110;
  assign T110 = acqNet_io_in_1_ready;
  assign io_clients_1_release_ready = T111;
  assign T111 = relNet_io_in_2_ready;
  assign io_clients_1_probe_bits_payload_p_type = T112;
  assign T112 = prbNet_io_out_2_bits_payload_p_type;
  assign io_clients_1_probe_bits_payload_addr = T113;
  assign T113 = prbNet_io_out_2_bits_payload_addr;
  assign io_clients_1_probe_bits_header_dst = T114;
  assign T114 = T115;
  assign T115 = prbNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_probe_bits_header_src = T116;
  assign T116 = prbNet_io_out_2_bits_header_src;
  assign io_clients_1_probe_valid = T117;
  assign T117 = prbNet_io_out_2_valid;
  assign io_clients_1_finish_ready = T118;
  assign T118 = ackNet_io_in_2_ready;
  assign io_clients_1_grant_bits_payload_g_type = T119;
  assign T119 = gntNet_io_out_2_bits_payload_g_type;
  assign io_clients_1_grant_bits_payload_uncached = T120;
  assign T120 = gntNet_io_out_2_bits_payload_uncached;
  assign io_clients_1_grant_bits_payload_manager_xact_id = T121;
  assign T121 = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign io_clients_1_grant_bits_payload_client_xact_id = T122;
  assign T122 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign io_clients_1_grant_bits_payload_data = T123;
  assign T123 = gntNet_io_out_2_bits_payload_data;
  assign io_clients_1_grant_bits_header_dst = T124;
  assign T124 = T125;
  assign T125 = gntNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_grant_bits_header_src = T126;
  assign T126 = gntNet_io_out_2_bits_header_src;
  assign io_clients_1_grant_valid = T127;
  assign T127 = gntNet_io_out_2_valid;
  assign io_clients_1_acquire_ready = T128;
  assign T128 = acqNet_io_in_2_ready;
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T67 ),
       .io_in_2_bits_header_src( T65 ),
       .io_in_2_bits_header_dst( T64 ),
       .io_in_2_bits_payload_addr( T63 ),
       .io_in_2_bits_payload_client_xact_id( T62 ),
       .io_in_2_bits_payload_data( T61 ),
       .io_in_2_bits_payload_uncached( T60 ),
       .io_in_2_bits_payload_a_type( T59 ),
       .io_in_2_bits_payload_subblock( T58 ),
       .io_in_1_ready( acqNet_io_in_1_ready ),
       .io_in_1_valid( T57 ),
       .io_in_1_bits_header_src( T55 ),
       .io_in_1_bits_header_dst( T54 ),
       .io_in_1_bits_payload_addr( T53 ),
       .io_in_1_bits_payload_client_xact_id( T52 ),
       .io_in_1_bits_payload_data( T51 ),
       .io_in_1_bits_payload_uncached( T50 ),
       .io_in_1_bits_payload_a_type( T49 ),
       .io_in_1_bits_payload_subblock( T48 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_uncached(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_subblock(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_uncached(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_subblock(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_uncached(  )
       //.io_out_1_bits_payload_a_type(  )
       //.io_out_1_bits_payload_subblock(  )
       .io_out_0_ready( T47 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( acqNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_uncached( acqNet_io_out_0_bits_payload_uncached ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_subblock( acqNet_io_out_0_bits_payload_subblock )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {5{$random}};
    assign acqNet.io_in_0_bits_payload_uncached = {1{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_subblock = {5{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T46 ),
       .io_in_2_bits_header_src( T44 ),
       .io_in_2_bits_header_dst( T43 ),
       .io_in_2_bits_payload_addr( T42 ),
       .io_in_2_bits_payload_client_xact_id( T41 ),
       .io_in_2_bits_payload_data( T40 ),
       .io_in_2_bits_payload_r_type( T39 ),
       .io_in_1_ready( relNet_io_in_1_ready ),
       .io_in_1_valid( T38 ),
       .io_in_1_bits_header_src( T36 ),
       .io_in_1_bits_header_dst( T35 ),
       .io_in_1_bits_payload_addr( T34 ),
       .io_in_1_bits_payload_client_xact_id( T33 ),
       .io_in_1_bits_payload_data( T32 ),
       .io_in_1_bits_payload_r_type( T31 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_r_type(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_r_type(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_r_type(  )
       .io_out_0_ready( T30 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( relNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {5{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr(  )
       //.io_in_2_bits_payload_p_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr(  )
       //.io_in_1_bits_payload_p_type(  )
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T29 ),
       .io_in_0_bits_header_src( T28 ),
       .io_in_0_bits_header_dst( T26 ),
       .io_in_0_bits_payload_addr( T25 ),
       .io_in_0_bits_payload_p_type( T24 ),
       .io_out_2_ready( T23 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr( prbNet_io_out_2_bits_payload_addr ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( T22 ),
       .io_out_1_valid( prbNet_io_out_1_valid ),
       .io_out_1_bits_header_src( prbNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( prbNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr( prbNet_io_out_1_bits_payload_addr ),
       .io_out_1_bits_payload_p_type( prbNet_io_out_1_bits_payload_p_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr(  )
       //.io_out_0_bits_payload_p_type(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_1_bits_header_src = {1{$random}};
    assign prbNet.io_in_1_bits_header_dst = {1{$random}};
    assign prbNet.io_in_1_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_1_bits_payload_p_type = {1{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_data(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_manager_xact_id(  )
       //.io_in_2_bits_payload_uncached(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_manager_xact_id(  )
       //.io_in_1_bits_payload_uncached(  )
       //.io_in_1_bits_payload_g_type(  )
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T21 ),
       .io_in_0_bits_header_src( T20 ),
       .io_in_0_bits_header_dst( T18 ),
       .io_in_0_bits_payload_data( T17 ),
       .io_in_0_bits_payload_client_xact_id( T16 ),
       .io_in_0_bits_payload_manager_xact_id( T15 ),
       .io_in_0_bits_payload_uncached( T14 ),
       .io_in_0_bits_payload_g_type( T13 ),
       .io_out_2_ready( T12 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_manager_xact_id( gntNet_io_out_2_bits_payload_manager_xact_id ),
       .io_out_2_bits_payload_uncached( gntNet_io_out_2_bits_payload_uncached ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_1_ready( T11 ),
       .io_out_1_valid( gntNet_io_out_1_valid ),
       .io_out_1_bits_header_src( gntNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( gntNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_data( gntNet_io_out_1_bits_payload_data ),
       .io_out_1_bits_payload_client_xact_id( gntNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_manager_xact_id( gntNet_io_out_1_bits_payload_manager_xact_id ),
       .io_out_1_bits_payload_uncached( gntNet_io_out_1_bits_payload_uncached ),
       .io_out_1_bits_payload_g_type( gntNet_io_out_1_bits_payload_g_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_data(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_manager_xact_id(  )
       //.io_out_0_bits_payload_uncached(  )
       //.io_out_0_bits_payload_g_type(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {5{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_manager_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_uncached = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_1_bits_header_src = {1{$random}};
    assign gntNet.io_in_1_bits_header_dst = {1{$random}};
    assign gntNet.io_in_1_bits_payload_data = {5{$random}};
    assign gntNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_manager_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_uncached = {1{$random}};
    assign gntNet.io_in_1_bits_payload_g_type = {1{$random}};
// synthesis translate_on
`endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( T8 ),
       .io_in_2_bits_header_dst( T7 ),
       .io_in_2_bits_payload_manager_xact_id( T6 ),
       .io_in_1_ready( ackNet_io_in_1_ready ),
       .io_in_1_valid( T5 ),
       .io_in_1_bits_header_src( T3 ),
       .io_in_1_bits_header_dst( T2 ),
       .io_in_1_bits_payload_manager_xact_id( T1 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_manager_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_manager_xact_id(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_manager_xact_id(  )
       .io_out_0_ready( T0 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_manager_xact_id( ackNet_io_out_0_bits_payload_manager_xact_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_manager_xact_id = {1{$random}};
// synthesis translate_on
`endif
endmodule

module VoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[1:0] io_inner_probe_bits_header_src
    //output[1:0] io_inner_probe_bits_header_dst
    //output[25:0] io_inner_probe_bits_payload_addr
    //output[1:0] io_inner_probe_bits_payload_p_type
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire[9:0] T1;
  wire[1:0] T2;
  wire T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  reg [3:0] xact_data_0;
  wire[3:0] T7;
  wire[3:0] T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[1:0] T12;
  reg [1:0] inner_data_cnt;
  wire[1:0] T104;
  wire[1:0] T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg  collect_inner_data;
  wire T105;
  wire T25;
  wire T26;
  wire T27;
  wire inner_data_done;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  reg [1:0] state;
  wire[1:0] T106;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire outer_data_done;
  wire T50;
  reg [1:0] outer_data_cnt;
  wire[1:0] T107;
  wire[1:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[3:0] T64;
  wire[1:0] T65;
  reg [3:0] xact_data_1;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[3:0] T74;
  reg [3:0] xact_data_2;
  wire[3:0] T75;
  wire[3:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  reg [3:0] xact_data_3;
  wire[3:0] T81;
  wire[3:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[4:0] T89;
  wire[25:0] T90;
  reg [25:0] xact_addr;
  wire[25:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[1:0] T97;
  wire T98;
  wire[3:0] T99;
  wire[1:0] T100;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T101;
  wire[3:0] T102;
  reg [1:0] xact_src;
  wire[1:0] T103;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    xact_data_0 = {1{$random}};
    inner_data_cnt = {1{$random}};
    collect_inner_data = {1{$random}};
    state = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    xact_addr = {1{$random}};
    xact_client_xact_id = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = io_inner_release_bits_payload_r_type == 3'h0;
  assign io_has_acquire_conflict = 1'h0;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = 1'h0;
  assign io_outer_acquire_bits_payload_subblock = T1;
  assign T1 = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T2;
  assign T2 = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T3;
  assign T3 = 1'h1;
  assign io_outer_acquire_bits_payload_data = T4;
  assign T4 = T5;
  assign T5 = T88 ? T74 : T6;
  assign T6 = T72 ? xact_data_1 : xact_data_0;
  assign T7 = T62 ? io_inner_release_bits_payload_data : T8;
  assign T8 = T9 ? io_inner_release_bits_payload_data : xact_data_0;
  assign T9 = T24 & T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = 1'h1 << T12;
  assign T12 = inner_data_cnt;
  assign T104 = reset ? 2'h0 : T13;
  assign T13 = T15 ? T14 : inner_data_cnt;
  assign T14 = inner_data_cnt + 2'h1;
  assign T15 = T23 & T16;
  assign T16 = T18 | T17;
  assign T17 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T18 = T20 | T19;
  assign T19 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T20 = T22 | T21;
  assign T21 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T22 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T23 = io_inner_release_ready & io_inner_release_valid;
  assign T24 = collect_inner_data & io_inner_release_valid;
  assign T105 = reset ? 1'h0 : T25;
  assign T25 = T36 ? T29 : T26;
  assign T26 = T27 ? 1'h0 : collect_inner_data;
  assign T27 = collect_inner_data & inner_data_done;
  assign inner_data_done = T15 & T28;
  assign T28 = inner_data_cnt == 2'h3;
  assign T29 = T31 | T30;
  assign T30 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T31 = T33 | T32;
  assign T32 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T33 = T35 | T34;
  assign T34 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T35 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T36 = T37 & io_inner_release_valid;
  assign T37 = 2'h0 == state;
  assign T106 = reset ? 2'h0 : T38;
  assign T38 = T60 ? 2'h0 : T39;
  assign T39 = T49 ? 2'h2 : T40;
  assign T40 = T36 ? T41 : state;
  assign T41 = T42 ? 2'h1 : 2'h2;
  assign T42 = T44 | T43;
  assign T43 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T46 = T48 | T47;
  assign T47 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T48 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T49 = T59 & outer_data_done;
  assign outer_data_done = T53 & T50;
  assign T50 = outer_data_cnt == 2'h3;
  assign T107 = reset ? 2'h0 : T51;
  assign T51 = T53 ? T52 : outer_data_cnt;
  assign T52 = outer_data_cnt + 2'h1;
  assign T53 = T58 & T54;
  assign T54 = io_outer_acquire_bits_payload_uncached ? T55 : 1'h0;
  assign T55 = T57 | T56;
  assign T56 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T57 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T58 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T59 = 2'h1 == state;
  assign T60 = T61 & io_inner_grant_ready;
  assign T61 = 2'h2 == state;
  assign T62 = T36 & T63;
  assign T63 = T64[1'h0:1'h0];
  assign T64 = 1'h1 << T65;
  assign T65 = 2'h0;
  assign T66 = T70 ? io_inner_release_bits_payload_data : T67;
  assign T67 = T68 ? io_inner_release_bits_payload_data : xact_data_1;
  assign T68 = T24 & T69;
  assign T69 = T11[1'h1:1'h1];
  assign T70 = T36 & T71;
  assign T71 = T64[1'h1:1'h1];
  assign T72 = T73[1'h0:1'h0];
  assign T73 = outer_data_cnt;
  assign T74 = T87 ? xact_data_3 : xact_data_2;
  assign T75 = T79 ? io_inner_release_bits_payload_data : T76;
  assign T76 = T77 ? io_inner_release_bits_payload_data : xact_data_2;
  assign T77 = T24 & T78;
  assign T78 = T11[2'h2:2'h2];
  assign T79 = T36 & T80;
  assign T80 = T64[2'h2:2'h2];
  assign T81 = T85 ? io_inner_release_bits_payload_data : T82;
  assign T82 = T83 ? io_inner_release_bits_payload_data : xact_data_3;
  assign T83 = T24 & T84;
  assign T84 = T11[2'h3:2'h3];
  assign T85 = T36 & T86;
  assign T86 = T64[2'h3:2'h3];
  assign T87 = T73[1'h0:1'h0];
  assign T88 = T73[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T89;
  assign T89 = 5'h0;
  assign io_outer_acquire_bits_payload_addr = T90;
  assign T90 = xact_addr;
  assign T91 = T36 ? io_inner_release_bits_payload_addr : xact_addr;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T92;
  assign T92 = T59 ? T93 : 1'h0;
  assign T93 = T95 | T94;
  assign T94 = outer_data_cnt < inner_data_cnt;
  assign T95 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T96;
  assign T96 = T37 ? 1'h1 : collect_inner_data;
//  assign io_inner_probe_bits_payload_p_type = {1{$random}};
//  assign io_inner_probe_bits_payload_addr = {1{$random}};
//  assign io_inner_probe_bits_header_dst = {1{$random}};
//  assign io_inner_probe_bits_header_src = {1{$random}};
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_finish_ready = 1'h0;
  assign io_inner_grant_bits_payload_g_type = T97;
  assign T97 = 2'h0;
  assign io_inner_grant_bits_payload_uncached = T98;
  assign T98 = 1'h0;
  assign io_inner_grant_bits_payload_manager_xact_id = T99;
  assign T99 = 4'h0;
  assign io_inner_grant_bits_payload_client_xact_id = T100;
  assign T100 = xact_client_xact_id;
  assign T101 = T36 ? io_inner_release_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T102;
  assign T102 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T103 = T36 ? io_inner_release_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T61;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(T62) begin
      xact_data_0 <= io_inner_release_bits_payload_data;
    end else if(T9) begin
      xact_data_0 <= io_inner_release_bits_payload_data;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T15) begin
      inner_data_cnt <= T14;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T36) begin
      collect_inner_data <= T29;
    end else if(T27) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T60) begin
      state <= 2'h0;
    end else if(T49) begin
      state <= 2'h2;
    end else if(T36) begin
      state <= T41;
    end
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T53) begin
      outer_data_cnt <= T52;
    end
    if(T70) begin
      xact_data_1 <= io_inner_release_bits_payload_data;
    end else if(T68) begin
      xact_data_1 <= io_inner_release_bits_payload_data;
    end
    if(T79) begin
      xact_data_2 <= io_inner_release_bits_payload_data;
    end else if(T77) begin
      xact_data_2 <= io_inner_release_bits_payload_data;
    end
    if(T85) begin
      xact_data_3 <= io_inner_release_bits_payload_data;
    end else if(T83) begin
      xact_data_3 <= io_inner_release_bits_payload_data;
    end
    if(T36) begin
      xact_addr <= io_inner_release_bits_payload_addr;
    end
    if(T36) begin
      xact_client_xact_id <= io_inner_release_bits_payload_client_xact_id;
    end
    if(T36) begin
      xact_src <= io_inner_release_bits_header_src;
    end
  end
endmodule

module AcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h1;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h1;
  assign outer_read_client_xact_id = 5'h1;
  assign outer_write_acq_client_xact_id = 5'h1;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h1;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h1;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module AcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h2;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h2;
  assign outer_read_client_xact_id = 5'h2;
  assign outer_write_acq_client_xact_id = 5'h2;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h2;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h2;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module AcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h3;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h3;
  assign outer_read_client_xact_id = 5'h3;
  assign outer_write_acq_client_xact_id = 5'h3;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h3;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h3;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module AcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h4;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h4;
  assign outer_read_client_xact_id = 5'h4;
  assign outer_write_acq_client_xact_id = 5'h4;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h4;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h4;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module AcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h5;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h5;
  assign outer_read_client_xact_id = 5'h5;
  assign outer_write_acq_client_xact_id = 5'h5;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h5;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h5;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module AcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h6;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h6;
  assign outer_read_client_xact_id = 5'h6;
  assign outer_write_acq_client_xact_id = 5'h6;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h6;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h6;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module AcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [3:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [9:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[3:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    //output[1:0] io_outer_acquire_bits_header_src
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[3:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[9:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [3:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output io_outer_finish_bits_payload_manager_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T224;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] myflag;
  wire[1:0] T21;
  wire T22;
  wire probe_self;
  wire T23;
  wire T24;
  wire T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire pending_outer_read;
  wire T28;
  wire[1:0] xact_a_type;
  reg [1:0] xact_a_type_;
  wire[1:0] T29;
  wire xact_uncached;
  reg  xact_uncached_;
  wire T30;
  wire pending_outer_write;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  release_count;
  wire T225;
  wire[1:0] T226;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T227;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T228;
  wire T42;
  wire[1:0] T229;
  wire T43;
  wire[1:0] T230;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire outer_data_done;
  wire T57;
  reg [1:0] outer_data_cnt;
  wire[1:0] T231;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[2:0] T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [25:0] xact_addr_;
  wire[25:0] T93;
  wire T94;
  wire T95;
  reg  collect_inner_data;
  wire T232;
  wire T96;
  wire T97;
  wire T98;
  wire inner_data_done;
  wire T99;
  reg [1:0] inner_data_cnt;
  wire[1:0] T233;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[9:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire[9:0] outer_write_rel_subblock;
  wire[9:0] outer_read_subblock;
  wire[9:0] outer_write_acq_subblock;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] outer_write_rel_a_type;
  wire[1:0] outer_read_a_type;
  wire[1:0] outer_write_acq_a_type;
  wire T121;
  wire T122;
  wire T123;
  wire outer_write_rel_uncached;
  wire outer_read_uncached;
  wire outer_write_acq_uncached;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_read_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T127;
  wire[3:0] T128;
  reg [3:0] xact_data_0;
  wire[3:0] T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg [3:0] xact_data_1;
  wire[3:0] T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire[3:0] T148;
  reg [3:0] xact_data_2;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  reg [3:0] xact_data_3;
  wire[3:0] T155;
  wire[3:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[4:0] T163;
  wire[4:0] T164;
  wire[4:0] T165;
  wire[4:0] outer_write_rel_client_xact_id;
  wire[4:0] outer_read_client_xact_id;
  wire[4:0] outer_write_acq_client_xact_id;
  wire[25:0] T166;
  wire[25:0] T167;
  wire[25:0] T168;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[25:0] T194;
  wire[1:0] T234;
  wire T235;
  wire T236;
  reg [1:0] probe_flags;
  wire[1:0] T237;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire[1:0] T215;
  reg [1:0] xact_client_xact_id_;
  wire[1:0] T216;
  wire[3:0] T217;
  reg [1:0] xact_src;
  wire[1:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type_ = {1{$random}};
    xact_uncached_ = {1{$random}};
    release_count = {1{$random}};
    outer_data_cnt = {1{$random}};
    xact_addr_ = {1{$random}};
    collect_inner_data = {1{$random}};
    inner_data_cnt = {1{$random}};
    xact_data_0 = {1{$random}};
    xact_data_1 = {1{$random}};
    xact_data_2 = {1{$random}};
    xact_data_3 = {1{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id_ = {1{$random}};
    xact_src = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_has_release_match = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T224 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T80 : T4;
  assign T4 = T78 ? T77 : T5;
  assign T5 = T75 ? T72 : T6;
  assign T6 = T70 ? T68 : T7;
  assign T7 = T34 ? T26 : T8;
  assign T8 = T24 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T14 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_uncached ? T13 : 1'h1;
  assign T13 = io_inner_acquire_bits_payload_a_type != 2'h1;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | myflag;
  assign myflag = probe_self ? 2'h0 : T21;
  assign T21 = 1'h1 << T22;
  assign T22 = io_inner_acquire_bits_header_src[1'h0:1'h0];
  assign probe_self = io_inner_acquire_bits_payload_uncached & T23;
  assign T23 = io_inner_acquire_bits_payload_a_type == 2'h0;
  assign T24 = T25 & io_inner_acquire_valid;
  assign T25 = 3'h0 == state;
  assign T26 = pending_outer_write ? 3'h3 : T27;
  assign T27 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_uncached ? T28 : 1'h1;
  assign T28 = xact_a_type != 2'h1;
  assign xact_a_type = xact_a_type_;
  assign T29 = T24 ? io_inner_acquire_bits_payload_a_type : xact_a_type_;
  assign xact_uncached = xact_uncached_;
  assign T30 = T24 ? io_inner_acquire_bits_payload_uncached : xact_uncached_;
  assign pending_outer_write = xact_uncached ? T31 : 1'h0;
  assign T31 = T33 | T32;
  assign T32 = 2'h2 == xact_a_type;
  assign T33 = 2'h1 == xact_a_type;
  assign T34 = T56 & T35;
  assign T35 = release_count == 1'h1;
  assign T225 = T226[1'h0:1'h0];
  assign T226 = reset ? 2'h0 : T36;
  assign T36 = T45 ? T230 : T37;
  assign T37 = T56 ? T229 : T38;
  assign T38 = T24 ? T39 : T227;
  assign T227 = {1'h0, release_count};
  assign T39 = T228 + T40;
  assign T40 = {1'h0, T41};
  assign T41 = probe_initial_flags[1'h1:1'h1];
  assign T228 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h0:1'h0];
  assign T229 = {1'h0, T43};
  assign T43 = release_count - 1'h1;
  assign T230 = {1'h0, T44};
  assign T44 = release_count - 1'h1;
  assign T45 = T54 & T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T49 | T48;
  assign T48 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T53 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T54 = T55 & io_inner_release_valid;
  assign T55 = 3'h1 == state;
  assign T56 = T66 & outer_data_done;
  assign outer_data_done = T60 & T57;
  assign T57 = outer_data_cnt == 2'h3;
  assign T231 = reset ? 2'h0 : T58;
  assign T58 = T60 ? T59 : outer_data_cnt;
  assign T59 = outer_data_cnt + 2'h1;
  assign T60 = T65 & T61;
  assign T61 = io_outer_acquire_bits_payload_uncached ? T62 : 1'h0;
  assign T62 = T64 | T63;
  assign T63 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T64 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T65 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T66 = T67 & io_outer_acquire_ready;
  assign T67 = T54 & T47;
  assign T68 = pending_outer_write ? 3'h3 : T69;
  assign T69 = pending_outer_read ? 3'h2 : 3'h4;
  assign T70 = T45 & T71;
  assign T71 = release_count == 1'h1;
  assign T72 = T73 ? 3'h5 : 3'h0;
  assign T73 = io_inner_grant_bits_payload_uncached | T74;
  assign T74 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T75 = T76 & io_outer_acquire_ready;
  assign T76 = 3'h2 == state;
  assign T77 = pending_outer_read ? 3'h2 : 3'h4;
  assign T78 = T79 & outer_data_done;
  assign T79 = 3'h3 == state;
  assign T80 = T81 ? 3'h5 : 3'h0;
  assign T81 = io_inner_grant_bits_payload_uncached | T82;
  assign T82 = io_inner_grant_bits_payload_g_type != 2'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_manager_xact_id == 4'h7;
  assign T88 = 3'h5 == state;
  assign T89 = T92 & T90;
  assign T90 = T91 ^ 1'h1;
  assign T91 = io_inner_release_bits_payload_r_type == 3'h0;
  assign T92 = xact_addr_ == io_inner_release_bits_payload_addr;
  assign T93 = T24 ? io_inner_acquire_bits_payload_addr : xact_addr_;
  assign io_has_acquire_conflict = T94;
  assign T94 = T112 & T95;
  assign T95 = collect_inner_data ^ 1'h1;
  assign T232 = reset ? 1'h0 : T96;
  assign T96 = T24 ? T108 : T97;
  assign T97 = T98 ? 1'h0 : collect_inner_data;
  assign T98 = collect_inner_data & inner_data_done;
  assign inner_data_done = T102 & T99;
  assign T99 = inner_data_cnt == 2'h3;
  assign T233 = reset ? 2'h0 : T100;
  assign T100 = T102 ? T101 : inner_data_cnt;
  assign T101 = inner_data_cnt + 2'h1;
  assign T102 = T107 & T103;
  assign T103 = io_inner_acquire_bits_payload_uncached ? T104 : 1'h0;
  assign T104 = T106 | T105;
  assign T105 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T106 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T107 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T108 = io_inner_acquire_bits_payload_uncached ? T109 : 1'h0;
  assign T109 = T111 | T110;
  assign T110 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T111 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T112 = T114 & T113;
  assign T113 = state != 3'h0;
  assign T114 = xact_addr_ == io_inner_acquire_bits_payload_addr;
//  assign io_outer_finish_bits_payload_manager_xact_id = {1{$random}};
//  assign io_outer_finish_bits_header_dst = {1{$random}};
//  assign io_outer_finish_bits_header_src = {1{$random}};
//  assign io_outer_finish_valid = {1{$random}};
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T115;
  assign T115 = T79 ? outer_write_acq_subblock : T116;
  assign T116 = T76 ? outer_read_subblock : T117;
  assign T117 = T67 ? outer_write_rel_subblock : outer_read_subblock;
  assign outer_write_rel_subblock = 10'h3;
  assign outer_read_subblock = 10'hf;
  assign outer_write_acq_subblock = 10'h3;
  assign io_outer_acquire_bits_payload_a_type = T118;
  assign T118 = T79 ? outer_write_acq_a_type : T119;
  assign T119 = T76 ? outer_read_a_type : T120;
  assign T120 = T67 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 2'h1;
  assign outer_read_a_type = 2'h0;
  assign outer_write_acq_a_type = 2'h1;
  assign io_outer_acquire_bits_payload_uncached = T121;
  assign T121 = T79 ? outer_write_acq_uncached : T122;
  assign T122 = T76 ? outer_read_uncached : T123;
  assign T123 = T67 ? outer_write_rel_uncached : outer_read_uncached;
  assign outer_write_rel_uncached = 1'h1;
  assign outer_read_uncached = 1'h1;
  assign outer_write_acq_uncached = 1'h1;
  assign io_outer_acquire_bits_payload_data = T124;
  assign T124 = T79 ? outer_write_acq_data : T125;
  assign T125 = T76 ? outer_read_data : T126;
  assign T126 = T67 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 4'h0;
  assign outer_write_acq_data = T127;
  assign T127 = T162 ? T148 : T128;
  assign T128 = T146 ? xact_data_1 : xact_data_0;
  assign T129 = T136 ? io_inner_acquire_bits_payload_data : T130;
  assign T130 = T131 ? io_inner_acquire_bits_payload_data : xact_data_0;
  assign T131 = T135 & T132;
  assign T132 = T133[1'h0:1'h0];
  assign T133 = 1'h1 << T134;
  assign T134 = inner_data_cnt;
  assign T135 = collect_inner_data & io_inner_acquire_valid;
  assign T136 = T24 & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = 2'h0;
  assign T140 = T144 ? io_inner_acquire_bits_payload_data : T141;
  assign T141 = T142 ? io_inner_acquire_bits_payload_data : xact_data_1;
  assign T142 = T135 & T143;
  assign T143 = T133[1'h1:1'h1];
  assign T144 = T24 & T145;
  assign T145 = T138[1'h1:1'h1];
  assign T146 = T147[1'h0:1'h0];
  assign T147 = outer_data_cnt;
  assign T148 = T161 ? xact_data_3 : xact_data_2;
  assign T149 = T153 ? io_inner_acquire_bits_payload_data : T150;
  assign T150 = T151 ? io_inner_acquire_bits_payload_data : xact_data_2;
  assign T151 = T135 & T152;
  assign T152 = T133[2'h2:2'h2];
  assign T153 = T24 & T154;
  assign T154 = T138[2'h2:2'h2];
  assign T155 = T159 ? io_inner_acquire_bits_payload_data : T156;
  assign T156 = T157 ? io_inner_acquire_bits_payload_data : xact_data_3;
  assign T157 = T135 & T158;
  assign T158 = T133[2'h3:2'h3];
  assign T159 = T24 & T160;
  assign T160 = T138[2'h3:2'h3];
  assign T161 = T147[1'h0:1'h0];
  assign T162 = T147[1'h1:1'h1];
  assign io_outer_acquire_bits_payload_client_xact_id = T163;
  assign T163 = T79 ? outer_write_acq_client_xact_id : T164;
  assign T164 = T76 ? outer_read_client_xact_id : T165;
  assign T165 = T67 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 5'h7;
  assign outer_read_client_xact_id = 5'h7;
  assign outer_write_acq_client_xact_id = 5'h7;
  assign io_outer_acquire_bits_payload_addr = T166;
  assign T166 = T79 ? outer_write_acq_addr : T167;
  assign T167 = T76 ? outer_read_addr : T168;
  assign T168 = T67 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr_;
  assign outer_read_addr = xact_addr_;
  assign outer_write_acq_addr = xact_addr_;
//  assign io_outer_acquire_bits_header_dst = {1{$random}};
//  assign io_outer_acquire_bits_header_src = {1{$random}};
  assign io_outer_acquire_valid = T169;
  assign T169 = T79 ? T171 : T170;
  assign T170 = T76 ? 1'h1 : T67;
  assign T171 = T173 | T172;
  assign T172 = outer_data_cnt < inner_data_cnt;
  assign T173 = collect_inner_data ^ 1'h1;
  assign io_inner_release_ready = T174;
  assign T174 = T55 ? T175 : 1'h0;
  assign T175 = T176 | io_outer_acquire_ready;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T179 | T178;
  assign T178 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T179 = T181 | T180;
  assign T180 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T181 = T183 | T182;
  assign T182 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T183 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign io_inner_probe_bits_payload_p_type = T184;
  assign T184 = T185;
  assign T185 = xact_uncached ? T188 : T186;
  assign T186 = T187 ? 2'h1 : 2'h0;
  assign T187 = xact_a_type == 2'h0;
  assign T188 = T193 ? 2'h2 : T189;
  assign T189 = T192 ? 2'h0 : T190;
  assign T190 = T191 ? 2'h0 : 2'h2;
  assign T191 = xact_a_type == 2'h2;
  assign T192 = xact_a_type == 2'h1;
  assign T193 = xact_a_type == 2'h0;
  assign io_inner_probe_bits_payload_addr = T194;
  assign T194 = xact_addr_;
  assign io_inner_probe_bits_header_dst = T234;
  assign T234 = {1'h0, T235};
  assign T235 = T236 == 1'h0;
  assign T236 = probe_flags[1'h0:1'h0];
  assign T237 = reset ? 2'h0 : T195;
  assign T195 = T200 ? T197 : T196;
  assign T196 = T24 ? probe_initial_flags : probe_flags;
  assign T197 = probe_flags & T198;
  assign T198 = ~ T199;
  assign T199 = 1'h1 << T235;
  assign T200 = T55 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T201;
  assign T201 = T55 ? T202 : 1'h0;
  assign T202 = probe_flags != 2'h0;
//  assign io_inner_finish_ready = {1{$random}};
  assign io_inner_grant_bits_payload_g_type = T203;
  assign T203 = T204;
  assign T204 = xact_uncached ? T207 : T205;
  assign T205 = T206 ? 2'h1 : 2'h2;
  assign T206 = xact_a_type == 2'h0;
  assign T207 = T212 ? 2'h0 : T208;
  assign T208 = T211 ? 2'h1 : T209;
  assign T209 = T210 ? 2'h2 : 2'h0;
  assign T210 = xact_a_type == 2'h2;
  assign T211 = xact_a_type == 2'h1;
  assign T212 = xact_a_type == 2'h0;
  assign io_inner_grant_bits_payload_uncached = T213;
  assign T213 = xact_uncached_;
  assign io_inner_grant_bits_payload_manager_xact_id = T214;
  assign T214 = 4'h7;
  assign io_inner_grant_bits_payload_client_xact_id = T215;
  assign T215 = xact_client_xact_id_;
  assign T216 = T24 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id_;
  assign io_inner_grant_bits_payload_data = T217;
  assign T217 = 4'h0;
  assign io_inner_grant_bits_header_dst = xact_src;
  assign T218 = T24 ? io_inner_acquire_bits_header_src : xact_src;
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T219;
  assign T219 = T220 ? 1'h1 : T84;
  assign T220 = T88 & T221;
  assign T221 = io_outer_grant_valid & T222;
  assign T222 = io_outer_grant_bits_payload_client_xact_id == 5'h7;
  assign io_inner_acquire_ready = T223;
  assign T223 = T25 ? 1'h1 : collect_inner_data;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T80;
    end else if(T78) begin
      state <= T77;
    end else if(T75) begin
      state <= T72;
    end else if(T70) begin
      state <= T68;
    end else if(T34) begin
      state <= T26;
    end else if(T24) begin
      state <= T9;
    end
    if(T24) begin
      xact_a_type_ <= io_inner_acquire_bits_payload_a_type;
    end
    if(T24) begin
      xact_uncached_ <= io_inner_acquire_bits_payload_uncached;
    end
    release_count <= T225;
    if(reset) begin
      outer_data_cnt <= 2'h0;
    end else if(T60) begin
      outer_data_cnt <= T59;
    end
    if(T24) begin
      xact_addr_ <= io_inner_acquire_bits_payload_addr;
    end
    if(reset) begin
      collect_inner_data <= 1'h0;
    end else if(T24) begin
      collect_inner_data <= T108;
    end else if(T98) begin
      collect_inner_data <= 1'h0;
    end
    if(reset) begin
      inner_data_cnt <= 2'h0;
    end else if(T102) begin
      inner_data_cnt <= T101;
    end
    if(T136) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end else if(T131) begin
      xact_data_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T144) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end else if(T142) begin
      xact_data_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T153) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end else if(T151) begin
      xact_data_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T159) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end else if(T157) begin
      xact_data_3 <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T200) begin
      probe_flags <= T197;
    end else if(T24) begin
      probe_flags <= probe_initial_flags;
    end
    if(T24) begin
      xact_client_xact_id_ <= io_inner_acquire_bits_payload_client_xact_id;
    end
    if(T24) begin
      xact_src <= io_inner_acquire_bits_header_src;
    end
  end
endmodule

module Arbiter_9(
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : T3;
  assign T3 = io_in_4_valid ? 3'h4 : T4;
  assign T4 = io_in_5_valid ? 3'h5 : T5;
  assign T5 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits = T6;
  assign T6 = T20 ? T14 : T7;
  assign T7 = T13 ? T11 : T8;
  assign T8 = T9 ? io_in_1_bits : io_in_0_bits;
  assign T9 = T10[1'h0:1'h0];
  assign T10 = chosen;
  assign T11 = T12 ? io_in_3_bits : io_in_2_bits;
  assign T12 = T10[1'h0:1'h0];
  assign T13 = T10[1'h1:1'h1];
  assign T14 = T19 ? T17 : T15;
  assign T15 = T16 ? io_in_5_bits : io_in_4_bits;
  assign T16 = T10[1'h0:1'h0];
  assign T17 = T18 ? io_in_7_bits : io_in_6_bits;
  assign T18 = T10[1'h0:1'h0];
  assign T19 = T10[1'h1:1'h1];
  assign T20 = T10[2'h2:2'h2];
  assign io_out_valid = T21;
  assign T21 = T34 ? T28 : T22;
  assign T22 = T27 ? T25 : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T10[1'h0:1'h0];
  assign T25 = T26 ? io_in_3_valid : io_in_2_valid;
  assign T26 = T10[1'h0:1'h0];
  assign T27 = T10[1'h1:1'h1];
  assign T28 = T33 ? T31 : T29;
  assign T29 = T30 ? io_in_5_valid : io_in_4_valid;
  assign T30 = T10[1'h0:1'h0];
  assign T31 = T32 ? io_in_7_valid : io_in_6_valid;
  assign T32 = T10[1'h0:1'h0];
  assign T33 = T10[1'h1:1'h1];
  assign T34 = T10[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T35;
  assign T35 = T36 & io_out_ready;
  assign T36 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = T39 ^ 1'h1;
  assign T39 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T40;
  assign T40 = T41 & io_out_ready;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T43 | io_in_2_valid;
  assign T43 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T44;
  assign T44 = T45 & io_out_ready;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 | io_in_3_valid;
  assign T47 = T48 | io_in_2_valid;
  assign T48 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T49;
  assign T49 = T50 & io_out_ready;
  assign T50 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_4_valid;
  assign T52 = T53 | io_in_3_valid;
  assign T53 = T54 | io_in_2_valid;
  assign T54 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T55;
  assign T55 = T56 & io_out_ready;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T58 | io_in_5_valid;
  assign T58 = T59 | io_in_4_valid;
  assign T59 = T60 | io_in_3_valid;
  assign T60 = T61 | io_in_2_valid;
  assign T61 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T62;
  assign T62 = T63 & io_out_ready;
  assign T63 = T64 ^ 1'h1;
  assign T64 = T65 | io_in_6_valid;
  assign T65 = T66 | io_in_5_valid;
  assign T66 = T67 | io_in_4_valid;
  assign T67 = T68 | io_in_3_valid;
  assign T68 = T69 | io_in_2_valid;
  assign T69 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_10(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [1:0] io_in_7_bits_payload_p_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [1:0] io_in_6_bits_payload_p_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [1:0] io_in_5_bits_payload_p_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire T9;
  wire[2:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire[25:0] T21;
  wire[25:0] T22;
  wire[25:0] T23;
  wire T24;
  wire[25:0] T25;
  wire T26;
  wire T27;
  wire[25:0] T28;
  wire[25:0] T29;
  wire T30;
  wire[25:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : T3;
  assign T3 = io_in_4_valid ? 3'h4 : T4;
  assign T4 = io_in_5_valid ? 3'h5 : T5;
  assign T5 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_p_type = T6;
  assign T6 = T20 ? T14 : T7;
  assign T7 = T13 ? T11 : T8;
  assign T8 = T9 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T9 = T10[1'h0:1'h0];
  assign T10 = chosen;
  assign T11 = T12 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T12 = T10[1'h0:1'h0];
  assign T13 = T10[1'h1:1'h1];
  assign T14 = T19 ? T17 : T15;
  assign T15 = T16 ? io_in_5_bits_payload_p_type : io_in_4_bits_payload_p_type;
  assign T16 = T10[1'h0:1'h0];
  assign T17 = T18 ? io_in_7_bits_payload_p_type : io_in_6_bits_payload_p_type;
  assign T18 = T10[1'h0:1'h0];
  assign T19 = T10[1'h1:1'h1];
  assign T20 = T10[2'h2:2'h2];
  assign io_out_bits_payload_addr = T21;
  assign T21 = T34 ? T28 : T22;
  assign T22 = T27 ? T25 : T23;
  assign T23 = T24 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T24 = T10[1'h0:1'h0];
  assign T25 = T26 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T26 = T10[1'h0:1'h0];
  assign T27 = T10[1'h1:1'h1];
  assign T28 = T33 ? T31 : T29;
  assign T29 = T30 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T30 = T10[1'h0:1'h0];
  assign T31 = T32 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T32 = T10[1'h0:1'h0];
  assign T33 = T10[1'h1:1'h1];
  assign T34 = T10[2'h2:2'h2];
  assign io_out_bits_header_dst = T35;
  assign T35 = T48 ? T42 : T36;
  assign T36 = T41 ? T39 : T37;
  assign T37 = T38 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T38 = T10[1'h0:1'h0];
  assign T39 = T40 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T40 = T10[1'h0:1'h0];
  assign T41 = T10[1'h1:1'h1];
  assign T42 = T47 ? T45 : T43;
  assign T43 = T44 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T44 = T10[1'h0:1'h0];
  assign T45 = T46 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T46 = T10[1'h0:1'h0];
  assign T47 = T10[1'h1:1'h1];
  assign T48 = T10[2'h2:2'h2];
  assign io_out_bits_header_src = T49;
  assign T49 = T62 ? T56 : T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T52 = T10[1'h0:1'h0];
  assign T53 = T54 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T54 = T10[1'h0:1'h0];
  assign T55 = T10[1'h1:1'h1];
  assign T56 = T61 ? T59 : T57;
  assign T57 = T58 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T58 = T10[1'h0:1'h0];
  assign T59 = T60 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T60 = T10[1'h0:1'h0];
  assign T61 = T10[1'h1:1'h1];
  assign T62 = T10[2'h2:2'h2];
  assign io_out_valid = T63;
  assign T63 = T76 ? T70 : T64;
  assign T64 = T69 ? T67 : T65;
  assign T65 = T66 ? io_in_1_valid : io_in_0_valid;
  assign T66 = T10[1'h0:1'h0];
  assign T67 = T68 ? io_in_3_valid : io_in_2_valid;
  assign T68 = T10[1'h0:1'h0];
  assign T69 = T10[1'h1:1'h1];
  assign T70 = T75 ? T73 : T71;
  assign T71 = T72 ? io_in_5_valid : io_in_4_valid;
  assign T72 = T10[1'h0:1'h0];
  assign T73 = T74 ? io_in_7_valid : io_in_6_valid;
  assign T74 = T10[1'h0:1'h0];
  assign T75 = T10[1'h1:1'h1];
  assign T76 = T10[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T77;
  assign T77 = T78 & io_out_ready;
  assign T78 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T79;
  assign T79 = T80 & io_out_ready;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T82;
  assign T82 = T83 & io_out_ready;
  assign T83 = T84 ^ 1'h1;
  assign T84 = T85 | io_in_2_valid;
  assign T85 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T86;
  assign T86 = T87 & io_out_ready;
  assign T87 = T88 ^ 1'h1;
  assign T88 = T89 | io_in_3_valid;
  assign T89 = T90 | io_in_2_valid;
  assign T90 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T91;
  assign T91 = T92 & io_out_ready;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T94 | io_in_4_valid;
  assign T94 = T95 | io_in_3_valid;
  assign T95 = T96 | io_in_2_valid;
  assign T96 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T97;
  assign T97 = T98 & io_out_ready;
  assign T98 = T99 ^ 1'h1;
  assign T99 = T100 | io_in_5_valid;
  assign T100 = T101 | io_in_4_valid;
  assign T101 = T102 | io_in_3_valid;
  assign T102 = T103 | io_in_2_valid;
  assign T103 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T104;
  assign T104 = T105 & io_out_ready;
  assign T105 = T106 ^ 1'h1;
  assign T106 = T107 | io_in_6_valid;
  assign T107 = T108 | io_in_5_valid;
  assign T108 = T109 | io_in_4_valid;
  assign T109 = T110 | io_in_3_valid;
  assign T110 = T111 | io_in_2_valid;
  assign T111 = io_in_0_valid | io_in_1_valid;
endmodule

module LockingArbiter_2(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [135:0] io_in_7_bits_payload_data,
    input [1:0] io_in_7_bits_payload_client_xact_id,
    input [3:0] io_in_7_bits_payload_manager_xact_id,
    input  io_in_7_bits_payload_uncached,
    input [1:0] io_in_7_bits_payload_g_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [135:0] io_in_6_bits_payload_data,
    input [1:0] io_in_6_bits_payload_client_xact_id,
    input [3:0] io_in_6_bits_payload_manager_xact_id,
    input  io_in_6_bits_payload_uncached,
    input [1:0] io_in_6_bits_payload_g_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [135:0] io_in_5_bits_payload_data,
    input [1:0] io_in_5_bits_payload_client_xact_id,
    input [3:0] io_in_5_bits_payload_manager_xact_id,
    input  io_in_5_bits_payload_uncached,
    input [1:0] io_in_5_bits_payload_g_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [135:0] io_in_4_bits_payload_data,
    input [1:0] io_in_4_bits_payload_client_xact_id,
    input [3:0] io_in_4_bits_payload_manager_xact_id,
    input  io_in_4_bits_payload_uncached,
    input [1:0] io_in_4_bits_payload_g_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [135:0] io_in_3_bits_payload_data,
    input [1:0] io_in_3_bits_payload_client_xact_id,
    input [3:0] io_in_3_bits_payload_manager_xact_id,
    input  io_in_3_bits_payload_uncached,
    input [1:0] io_in_3_bits_payload_g_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [135:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_manager_xact_id,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [135:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_manager_xact_id,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [135:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_manager_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[135:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_manager_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  reg [2:0] lockIdx;
  wire[2:0] T205;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  locked;
  wire T206;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  reg [1:0] R38;
  wire[1:0] T207;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire[2:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire[3:0] T76;
  wire[3:0] T77;
  wire T78;
  wire[3:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[1:0] T87;
  wire T88;
  wire T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire T92;
  wire[1:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire[135:0] T97;
  wire[135:0] T98;
  wire[135:0] T99;
  wire T100;
  wire[135:0] T101;
  wire T102;
  wire T103;
  wire[135:0] T104;
  wire[135:0] T105;
  wire T106;
  wire[135:0] T107;
  wire T108;
  wire T109;
  wire T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] T113;
  wire T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire T120;
  wire[1:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire T128;
  wire[1:0] T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R38 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid ? 3'h0 : T1;
  assign T1 = io_in_1_valid ? 3'h1 : T2;
  assign T2 = io_in_2_valid ? 3'h2 : T3;
  assign T3 = io_in_3_valid ? 3'h3 : T4;
  assign T4 = io_in_4_valid ? 3'h4 : T5;
  assign T5 = io_in_5_valid ? 3'h5 : T6;
  assign T6 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T205 = reset ? 3'h7 : T7;
  assign T7 = T22 ? T8 : lockIdx;
  assign T8 = T21 ? 3'h0 : T9;
  assign T9 = T20 ? 3'h1 : T10;
  assign T10 = T19 ? 3'h2 : T11;
  assign T11 = T18 ? 3'h3 : T12;
  assign T12 = T17 ? 3'h4 : T13;
  assign T13 = T16 ? 3'h5 : T14;
  assign T14 = T15 ? 3'h6 : 3'h7;
  assign T15 = io_in_6_ready & io_in_6_valid;
  assign T16 = io_in_5_ready & io_in_5_valid;
  assign T17 = io_in_4_ready & io_in_4_valid;
  assign T18 = io_in_3_ready & io_in_3_valid;
  assign T19 = io_in_2_ready & io_in_2_valid;
  assign T20 = io_in_1_ready & io_in_1_valid;
  assign T21 = io_in_0_ready & io_in_0_valid;
  assign T22 = T24 & T23;
  assign T23 = locked ^ 1'h1;
  assign T24 = T32 & T25;
  assign T25 = io_out_bits_payload_uncached ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 2'h2 == io_out_bits_payload_g_type;
  assign T28 = 2'h1 == io_out_bits_payload_g_type;
  assign T29 = T31 | T30;
  assign T30 = 2'h2 == io_out_bits_payload_g_type;
  assign T31 = 2'h0 == io_out_bits_payload_g_type;
  assign T32 = io_out_ready & io_out_valid;
  assign T206 = reset ? 1'h0 : T33;
  assign T33 = T35 ? 1'h0 : T34;
  assign T34 = T22 ? 1'h1 : locked;
  assign T35 = T32 & T36;
  assign T36 = T37 == 2'h0;
  assign T37 = R38 + 2'h1;
  assign T207 = reset ? 2'h0 : T39;
  assign T39 = T24 ? T37 : R38;
  assign io_out_bits_payload_g_type = T40;
  assign T40 = T54 ? T48 : T41;
  assign T41 = T47 ? T45 : T42;
  assign T42 = T43 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T43 = T44[1'h0:1'h0];
  assign T44 = chosen;
  assign T45 = T46 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T46 = T44[1'h0:1'h0];
  assign T47 = T44[1'h1:1'h1];
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_5_bits_payload_g_type : io_in_4_bits_payload_g_type;
  assign T50 = T44[1'h0:1'h0];
  assign T51 = T52 ? io_in_7_bits_payload_g_type : io_in_6_bits_payload_g_type;
  assign T52 = T44[1'h0:1'h0];
  assign T53 = T44[1'h1:1'h1];
  assign T54 = T44[2'h2:2'h2];
  assign io_out_bits_payload_uncached = T55;
  assign T55 = T68 ? T62 : T56;
  assign T56 = T61 ? T59 : T57;
  assign T57 = T58 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T58 = T44[1'h0:1'h0];
  assign T59 = T60 ? io_in_3_bits_payload_uncached : io_in_2_bits_payload_uncached;
  assign T60 = T44[1'h0:1'h0];
  assign T61 = T44[1'h1:1'h1];
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_5_bits_payload_uncached : io_in_4_bits_payload_uncached;
  assign T64 = T44[1'h0:1'h0];
  assign T65 = T66 ? io_in_7_bits_payload_uncached : io_in_6_bits_payload_uncached;
  assign T66 = T44[1'h0:1'h0];
  assign T67 = T44[1'h1:1'h1];
  assign T68 = T44[2'h2:2'h2];
  assign io_out_bits_payload_manager_xact_id = T69;
  assign T69 = T82 ? T76 : T70;
  assign T70 = T75 ? T73 : T71;
  assign T71 = T72 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T72 = T44[1'h0:1'h0];
  assign T73 = T74 ? io_in_3_bits_payload_manager_xact_id : io_in_2_bits_payload_manager_xact_id;
  assign T74 = T44[1'h0:1'h0];
  assign T75 = T44[1'h1:1'h1];
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_5_bits_payload_manager_xact_id : io_in_4_bits_payload_manager_xact_id;
  assign T78 = T44[1'h0:1'h0];
  assign T79 = T80 ? io_in_7_bits_payload_manager_xact_id : io_in_6_bits_payload_manager_xact_id;
  assign T80 = T44[1'h0:1'h0];
  assign T81 = T44[1'h1:1'h1];
  assign T82 = T44[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T83;
  assign T83 = T96 ? T90 : T84;
  assign T84 = T89 ? T87 : T85;
  assign T85 = T86 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T86 = T44[1'h0:1'h0];
  assign T87 = T88 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T88 = T44[1'h0:1'h0];
  assign T89 = T44[1'h1:1'h1];
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T92 = T44[1'h0:1'h0];
  assign T93 = T94 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T94 = T44[1'h0:1'h0];
  assign T95 = T44[1'h1:1'h1];
  assign T96 = T44[2'h2:2'h2];
  assign io_out_bits_payload_data = T97;
  assign T97 = T110 ? T104 : T98;
  assign T98 = T103 ? T101 : T99;
  assign T99 = T100 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T100 = T44[1'h0:1'h0];
  assign T101 = T102 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T102 = T44[1'h0:1'h0];
  assign T103 = T44[1'h1:1'h1];
  assign T104 = T109 ? T107 : T105;
  assign T105 = T106 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T106 = T44[1'h0:1'h0];
  assign T107 = T108 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T108 = T44[1'h0:1'h0];
  assign T109 = T44[1'h1:1'h1];
  assign T110 = T44[2'h2:2'h2];
  assign io_out_bits_header_dst = T111;
  assign T111 = T124 ? T118 : T112;
  assign T112 = T117 ? T115 : T113;
  assign T113 = T114 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T114 = T44[1'h0:1'h0];
  assign T115 = T116 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T116 = T44[1'h0:1'h0];
  assign T117 = T44[1'h1:1'h1];
  assign T118 = T123 ? T121 : T119;
  assign T119 = T120 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T120 = T44[1'h0:1'h0];
  assign T121 = T122 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T122 = T44[1'h0:1'h0];
  assign T123 = T44[1'h1:1'h1];
  assign T124 = T44[2'h2:2'h2];
  assign io_out_bits_header_src = T125;
  assign T125 = T138 ? T132 : T126;
  assign T126 = T131 ? T129 : T127;
  assign T127 = T128 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T128 = T44[1'h0:1'h0];
  assign T129 = T130 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T130 = T44[1'h0:1'h0];
  assign T131 = T44[1'h1:1'h1];
  assign T132 = T137 ? T135 : T133;
  assign T133 = T134 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T134 = T44[1'h0:1'h0];
  assign T135 = T136 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T136 = T44[1'h0:1'h0];
  assign T137 = T44[1'h1:1'h1];
  assign T138 = T44[2'h2:2'h2];
  assign io_out_valid = T139;
  assign T139 = T152 ? T146 : T140;
  assign T140 = T145 ? T143 : T141;
  assign T141 = T142 ? io_in_1_valid : io_in_0_valid;
  assign T142 = T44[1'h0:1'h0];
  assign T143 = T144 ? io_in_3_valid : io_in_2_valid;
  assign T144 = T44[1'h0:1'h0];
  assign T145 = T44[1'h1:1'h1];
  assign T146 = T151 ? T149 : T147;
  assign T147 = T148 ? io_in_5_valid : io_in_4_valid;
  assign T148 = T44[1'h0:1'h0];
  assign T149 = T150 ? io_in_7_valid : io_in_6_valid;
  assign T150 = T44[1'h0:1'h0];
  assign T151 = T44[1'h1:1'h1];
  assign T152 = T44[2'h2:2'h2];
  assign io_in_0_ready = T153;
  assign T153 = T154 & io_out_ready;
  assign T154 = locked ? T155 : 1'h1;
  assign T155 = lockIdx == 3'h0;
  assign io_in_1_ready = T156;
  assign T156 = T157 & io_out_ready;
  assign T157 = locked ? T159 : T158;
  assign T158 = io_in_0_valid ^ 1'h1;
  assign T159 = lockIdx == 3'h1;
  assign io_in_2_ready = T160;
  assign T160 = T161 & io_out_ready;
  assign T161 = locked ? T164 : T162;
  assign T162 = T163 ^ 1'h1;
  assign T163 = io_in_0_valid | io_in_1_valid;
  assign T164 = lockIdx == 3'h2;
  assign io_in_3_ready = T165;
  assign T165 = T166 & io_out_ready;
  assign T166 = locked ? T170 : T167;
  assign T167 = T168 ^ 1'h1;
  assign T168 = T169 | io_in_2_valid;
  assign T169 = io_in_0_valid | io_in_1_valid;
  assign T170 = lockIdx == 3'h3;
  assign io_in_4_ready = T171;
  assign T171 = T172 & io_out_ready;
  assign T172 = locked ? T177 : T173;
  assign T173 = T174 ^ 1'h1;
  assign T174 = T175 | io_in_3_valid;
  assign T175 = T176 | io_in_2_valid;
  assign T176 = io_in_0_valid | io_in_1_valid;
  assign T177 = lockIdx == 3'h4;
  assign io_in_5_ready = T178;
  assign T178 = T179 & io_out_ready;
  assign T179 = locked ? T185 : T180;
  assign T180 = T181 ^ 1'h1;
  assign T181 = T182 | io_in_4_valid;
  assign T182 = T183 | io_in_3_valid;
  assign T183 = T184 | io_in_2_valid;
  assign T184 = io_in_0_valid | io_in_1_valid;
  assign T185 = lockIdx == 3'h5;
  assign io_in_6_ready = T186;
  assign T186 = T187 & io_out_ready;
  assign T187 = locked ? T194 : T188;
  assign T188 = T189 ^ 1'h1;
  assign T189 = T190 | io_in_5_valid;
  assign T190 = T191 | io_in_4_valid;
  assign T191 = T192 | io_in_3_valid;
  assign T192 = T193 | io_in_2_valid;
  assign T193 = io_in_0_valid | io_in_1_valid;
  assign T194 = lockIdx == 3'h6;
  assign io_in_7_ready = T195;
  assign T195 = T196 & io_out_ready;
  assign T196 = locked ? T204 : T197;
  assign T197 = T198 ^ 1'h1;
  assign T198 = T199 | io_in_6_valid;
  assign T199 = T200 | io_in_5_valid;
  assign T200 = T201 | io_in_4_valid;
  assign T201 = T202 | io_in_3_valid;
  assign T202 = T203 | io_in_2_valid;
  assign T203 = io_in_0_valid | io_in_1_valid;
  assign T204 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 3'h7;
    end else if(T22) begin
      lockIdx <= T8;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T35) begin
      locked <= 1'h0;
    end else if(T22) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R38 <= 2'h0;
    end else if(T24) begin
      R38 <= T37;
    end
  end
endmodule

module LockingRRArbiter_14(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [4:0] io_in_7_bits_payload_client_xact_id,
    input [3:0] io_in_7_bits_payload_data,
    input  io_in_7_bits_payload_uncached,
    input [1:0] io_in_7_bits_payload_a_type,
    input [9:0] io_in_7_bits_payload_subblock,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [4:0] io_in_6_bits_payload_client_xact_id,
    input [3:0] io_in_6_bits_payload_data,
    input  io_in_6_bits_payload_uncached,
    input [1:0] io_in_6_bits_payload_a_type,
    input [9:0] io_in_6_bits_payload_subblock,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [4:0] io_in_5_bits_payload_client_xact_id,
    input [3:0] io_in_5_bits_payload_data,
    input  io_in_5_bits_payload_uncached,
    input [1:0] io_in_5_bits_payload_a_type,
    input [9:0] io_in_5_bits_payload_subblock,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [4:0] io_in_4_bits_payload_client_xact_id,
    input [3:0] io_in_4_bits_payload_data,
    input  io_in_4_bits_payload_uncached,
    input [1:0] io_in_4_bits_payload_a_type,
    input [9:0] io_in_4_bits_payload_subblock,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [4:0] io_in_3_bits_payload_client_xact_id,
    input [3:0] io_in_3_bits_payload_data,
    input  io_in_3_bits_payload_uncached,
    input [1:0] io_in_3_bits_payload_a_type,
    input [9:0] io_in_3_bits_payload_subblock,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [4:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_uncached,
    input [1:0] io_in_2_bits_payload_a_type,
    input [9:0] io_in_2_bits_payload_subblock,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [4:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_uncached,
    input [1:0] io_in_1_bits_payload_a_type,
    input [9:0] io_in_1_bits_payload_subblock,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [4:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_a_type,
    input [9:0] io_in_0_bits_payload_subblock,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[4:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_data,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_a_type,
    output[9:0] io_out_bits_payload_subblock,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg [2:0] last_grant;
  wire[2:0] T370;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] lockIdx;
  wire[2:0] T371;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  reg  locked;
  wire T372;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  reg [1:0] R58;
  wire[1:0] T373;
  wire[1:0] T59;
  wire[9:0] T60;
  wire[9:0] T61;
  wire[9:0] T62;
  wire T63;
  wire[2:0] T64;
  wire[9:0] T65;
  wire T66;
  wire T67;
  wire[9:0] T68;
  wire[9:0] T69;
  wire T70;
  wire[9:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire T78;
  wire[1:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire[1:0] T83;
  wire T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[3:0] T103;
  wire[3:0] T104;
  wire[3:0] T105;
  wire T106;
  wire[3:0] T107;
  wire T108;
  wire T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire T112;
  wire[3:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[4:0] T117;
  wire[4:0] T118;
  wire[4:0] T119;
  wire T120;
  wire[4:0] T121;
  wire T122;
  wire T123;
  wire[4:0] T124;
  wire[4:0] T125;
  wire T126;
  wire[4:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[25:0] T131;
  wire[25:0] T132;
  wire[25:0] T133;
  wire T134;
  wire[25:0] T135;
  wire T136;
  wire T137;
  wire[25:0] T138;
  wire[25:0] T139;
  wire T140;
  wire[25:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[1:0] T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire T148;
  wire[1:0] T149;
  wire T150;
  wire T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[1:0] T163;
  wire T164;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire T168;
  wire[1:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R58 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T28 ? 3'h1 : T1;
  assign T1 = T26 ? 3'h2 : T2;
  assign T2 = T24 ? 3'h3 : T3;
  assign T3 = T22 ? 3'h4 : T4;
  assign T4 = T20 ? 3'h5 : T5;
  assign T5 = T18 ? 3'h6 : T6;
  assign T6 = T14 ? 3'h7 : T7;
  assign T7 = io_in_0_valid ? 3'h0 : T8;
  assign T8 = io_in_1_valid ? 3'h1 : T9;
  assign T9 = io_in_2_valid ? 3'h2 : T10;
  assign T10 = io_in_3_valid ? 3'h3 : T11;
  assign T11 = io_in_4_valid ? 3'h4 : T12;
  assign T12 = io_in_5_valid ? 3'h5 : T13;
  assign T13 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T14 = io_in_7_valid & T15;
  assign T15 = last_grant < 3'h7;
  assign T370 = reset ? 3'h0 : T16;
  assign T16 = T17 ? chosen : last_grant;
  assign T17 = io_out_ready & io_out_valid;
  assign T18 = io_in_6_valid & T19;
  assign T19 = last_grant < 3'h6;
  assign T20 = io_in_5_valid & T21;
  assign T21 = last_grant < 3'h5;
  assign T22 = io_in_4_valid & T23;
  assign T23 = last_grant < 3'h4;
  assign T24 = io_in_3_valid & T25;
  assign T25 = last_grant < 3'h3;
  assign T26 = io_in_2_valid & T27;
  assign T27 = last_grant < 3'h2;
  assign T28 = io_in_1_valid & T29;
  assign T29 = last_grant < 3'h1;
  assign T371 = reset ? 3'h7 : T30;
  assign T30 = T45 ? T31 : lockIdx;
  assign T31 = T44 ? 3'h0 : T32;
  assign T32 = T43 ? 3'h1 : T33;
  assign T33 = T42 ? 3'h2 : T34;
  assign T34 = T41 ? 3'h3 : T35;
  assign T35 = T40 ? 3'h4 : T36;
  assign T36 = T39 ? 3'h5 : T37;
  assign T37 = T38 ? 3'h6 : 3'h7;
  assign T38 = io_in_6_ready & io_in_6_valid;
  assign T39 = io_in_5_ready & io_in_5_valid;
  assign T40 = io_in_4_ready & io_in_4_valid;
  assign T41 = io_in_3_ready & io_in_3_valid;
  assign T42 = io_in_2_ready & io_in_2_valid;
  assign T43 = io_in_1_ready & io_in_1_valid;
  assign T44 = io_in_0_ready & io_in_0_valid;
  assign T45 = T47 & T46;
  assign T46 = locked ^ 1'h1;
  assign T47 = T52 & T48;
  assign T48 = io_out_bits_payload_uncached ? T49 : 1'h0;
  assign T49 = T51 | T50;
  assign T50 = 2'h2 == io_out_bits_payload_a_type;
  assign T51 = 2'h1 == io_out_bits_payload_a_type;
  assign T52 = io_out_ready & io_out_valid;
  assign T372 = reset ? 1'h0 : T53;
  assign T53 = T55 ? 1'h0 : T54;
  assign T54 = T45 ? 1'h1 : locked;
  assign T55 = T52 & T56;
  assign T56 = T57 == 2'h0;
  assign T57 = R58 + 2'h1;
  assign T373 = reset ? 2'h0 : T59;
  assign T59 = T47 ? T57 : R58;
  assign io_out_bits_payload_subblock = T60;
  assign T60 = T74 ? T68 : T61;
  assign T61 = T67 ? T65 : T62;
  assign T62 = T63 ? io_in_1_bits_payload_subblock : io_in_0_bits_payload_subblock;
  assign T63 = T64[1'h0:1'h0];
  assign T64 = chosen;
  assign T65 = T66 ? io_in_3_bits_payload_subblock : io_in_2_bits_payload_subblock;
  assign T66 = T64[1'h0:1'h0];
  assign T67 = T64[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_payload_subblock : io_in_4_bits_payload_subblock;
  assign T70 = T64[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_payload_subblock : io_in_6_bits_payload_subblock;
  assign T72 = T64[1'h0:1'h0];
  assign T73 = T64[1'h1:1'h1];
  assign T74 = T64[2'h2:2'h2];
  assign io_out_bits_payload_a_type = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T78 = T64[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T80 = T64[1'h0:1'h0];
  assign T81 = T64[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_bits_payload_a_type : io_in_4_bits_payload_a_type;
  assign T84 = T64[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_bits_payload_a_type : io_in_6_bits_payload_a_type;
  assign T86 = T64[1'h0:1'h0];
  assign T87 = T64[1'h1:1'h1];
  assign T88 = T64[2'h2:2'h2];
  assign io_out_bits_payload_uncached = T89;
  assign T89 = T102 ? T96 : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_payload_uncached : io_in_0_bits_payload_uncached;
  assign T92 = T64[1'h0:1'h0];
  assign T93 = T94 ? io_in_3_bits_payload_uncached : io_in_2_bits_payload_uncached;
  assign T94 = T64[1'h0:1'h0];
  assign T95 = T64[1'h1:1'h1];
  assign T96 = T101 ? T99 : T97;
  assign T97 = T98 ? io_in_5_bits_payload_uncached : io_in_4_bits_payload_uncached;
  assign T98 = T64[1'h0:1'h0];
  assign T99 = T100 ? io_in_7_bits_payload_uncached : io_in_6_bits_payload_uncached;
  assign T100 = T64[1'h0:1'h0];
  assign T101 = T64[1'h1:1'h1];
  assign T102 = T64[2'h2:2'h2];
  assign io_out_bits_payload_data = T103;
  assign T103 = T116 ? T110 : T104;
  assign T104 = T109 ? T107 : T105;
  assign T105 = T106 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T106 = T64[1'h0:1'h0];
  assign T107 = T108 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T108 = T64[1'h0:1'h0];
  assign T109 = T64[1'h1:1'h1];
  assign T110 = T115 ? T113 : T111;
  assign T111 = T112 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T112 = T64[1'h0:1'h0];
  assign T113 = T114 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T114 = T64[1'h0:1'h0];
  assign T115 = T64[1'h1:1'h1];
  assign T116 = T64[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T117;
  assign T117 = T130 ? T124 : T118;
  assign T118 = T123 ? T121 : T119;
  assign T119 = T120 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T120 = T64[1'h0:1'h0];
  assign T121 = T122 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T122 = T64[1'h0:1'h0];
  assign T123 = T64[1'h1:1'h1];
  assign T124 = T129 ? T127 : T125;
  assign T125 = T126 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T126 = T64[1'h0:1'h0];
  assign T127 = T128 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T128 = T64[1'h0:1'h0];
  assign T129 = T64[1'h1:1'h1];
  assign T130 = T64[2'h2:2'h2];
  assign io_out_bits_payload_addr = T131;
  assign T131 = T144 ? T138 : T132;
  assign T132 = T137 ? T135 : T133;
  assign T133 = T134 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T134 = T64[1'h0:1'h0];
  assign T135 = T136 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T136 = T64[1'h0:1'h0];
  assign T137 = T64[1'h1:1'h1];
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T140 = T64[1'h0:1'h0];
  assign T141 = T142 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T142 = T64[1'h0:1'h0];
  assign T143 = T64[1'h1:1'h1];
  assign T144 = T64[2'h2:2'h2];
  assign io_out_bits_header_dst = T145;
  assign T145 = T158 ? T152 : T146;
  assign T146 = T151 ? T149 : T147;
  assign T147 = T148 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T148 = T64[1'h0:1'h0];
  assign T149 = T150 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T150 = T64[1'h0:1'h0];
  assign T151 = T64[1'h1:1'h1];
  assign T152 = T157 ? T155 : T153;
  assign T153 = T154 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T154 = T64[1'h0:1'h0];
  assign T155 = T156 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T156 = T64[1'h0:1'h0];
  assign T157 = T64[1'h1:1'h1];
  assign T158 = T64[2'h2:2'h2];
  assign io_out_bits_header_src = T159;
  assign T159 = T172 ? T166 : T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T162 = T64[1'h0:1'h0];
  assign T163 = T164 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T164 = T64[1'h0:1'h0];
  assign T165 = T64[1'h1:1'h1];
  assign T166 = T171 ? T169 : T167;
  assign T167 = T168 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T168 = T64[1'h0:1'h0];
  assign T169 = T170 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T170 = T64[1'h0:1'h0];
  assign T171 = T64[1'h1:1'h1];
  assign T172 = T64[2'h2:2'h2];
  assign io_out_valid = T173;
  assign T173 = T186 ? T180 : T174;
  assign T174 = T179 ? T177 : T175;
  assign T175 = T176 ? io_in_1_valid : io_in_0_valid;
  assign T176 = T64[1'h0:1'h0];
  assign T177 = T178 ? io_in_3_valid : io_in_2_valid;
  assign T178 = T64[1'h0:1'h0];
  assign T179 = T64[1'h1:1'h1];
  assign T180 = T185 ? T183 : T181;
  assign T181 = T182 ? io_in_5_valid : io_in_4_valid;
  assign T182 = T64[1'h0:1'h0];
  assign T183 = T184 ? io_in_7_valid : io_in_6_valid;
  assign T184 = T64[1'h0:1'h0];
  assign T185 = T64[1'h1:1'h1];
  assign T186 = T64[2'h2:2'h2];
  assign io_in_0_ready = T187;
  assign T187 = T188 & io_out_ready;
  assign T188 = locked ? T215 : T189;
  assign T189 = T214 | T190;
  assign T190 = T191 ^ 1'h1;
  assign T191 = T194 | T192;
  assign T192 = io_in_7_valid & T193;
  assign T193 = last_grant < 3'h7;
  assign T194 = T197 | T195;
  assign T195 = io_in_6_valid & T196;
  assign T196 = last_grant < 3'h6;
  assign T197 = T200 | T198;
  assign T198 = io_in_5_valid & T199;
  assign T199 = last_grant < 3'h5;
  assign T200 = T203 | T201;
  assign T201 = io_in_4_valid & T202;
  assign T202 = last_grant < 3'h4;
  assign T203 = T206 | T204;
  assign T204 = io_in_3_valid & T205;
  assign T205 = last_grant < 3'h3;
  assign T206 = T209 | T207;
  assign T207 = io_in_2_valid & T208;
  assign T208 = last_grant < 3'h2;
  assign T209 = T212 | T210;
  assign T210 = io_in_1_valid & T211;
  assign T211 = last_grant < 3'h1;
  assign T212 = io_in_0_valid & T213;
  assign T213 = last_grant < 3'h0;
  assign T214 = last_grant < 3'h0;
  assign T215 = lockIdx == 3'h0;
  assign io_in_1_ready = T216;
  assign T216 = T217 & io_out_ready;
  assign T217 = locked ? T231 : T218;
  assign T218 = T228 | T219;
  assign T219 = T220 ^ 1'h1;
  assign T220 = T221 | io_in_0_valid;
  assign T221 = T222 | T192;
  assign T222 = T223 | T195;
  assign T223 = T224 | T198;
  assign T224 = T225 | T201;
  assign T225 = T226 | T204;
  assign T226 = T227 | T207;
  assign T227 = T212 | T210;
  assign T228 = T230 & T229;
  assign T229 = last_grant < 3'h1;
  assign T230 = T212 ^ 1'h1;
  assign T231 = lockIdx == 3'h1;
  assign io_in_2_ready = T232;
  assign T232 = T233 & io_out_ready;
  assign T233 = locked ? T249 : T234;
  assign T234 = T245 | T235;
  assign T235 = T236 ^ 1'h1;
  assign T236 = T237 | io_in_1_valid;
  assign T237 = T238 | io_in_0_valid;
  assign T238 = T239 | T192;
  assign T239 = T240 | T195;
  assign T240 = T241 | T198;
  assign T241 = T242 | T201;
  assign T242 = T243 | T204;
  assign T243 = T244 | T207;
  assign T244 = T212 | T210;
  assign T245 = T247 & T246;
  assign T246 = last_grant < 3'h2;
  assign T247 = T248 ^ 1'h1;
  assign T248 = T212 | T210;
  assign T249 = lockIdx == 3'h2;
  assign io_in_3_ready = T250;
  assign T250 = T251 & io_out_ready;
  assign T251 = locked ? T269 : T252;
  assign T252 = T264 | T253;
  assign T253 = T254 ^ 1'h1;
  assign T254 = T255 | io_in_2_valid;
  assign T255 = T256 | io_in_1_valid;
  assign T256 = T257 | io_in_0_valid;
  assign T257 = T258 | T192;
  assign T258 = T259 | T195;
  assign T259 = T260 | T198;
  assign T260 = T261 | T201;
  assign T261 = T262 | T204;
  assign T262 = T263 | T207;
  assign T263 = T212 | T210;
  assign T264 = T266 & T265;
  assign T265 = last_grant < 3'h3;
  assign T266 = T267 ^ 1'h1;
  assign T267 = T268 | T207;
  assign T268 = T212 | T210;
  assign T269 = lockIdx == 3'h3;
  assign io_in_4_ready = T270;
  assign T270 = T271 & io_out_ready;
  assign T271 = locked ? T291 : T272;
  assign T272 = T285 | T273;
  assign T273 = T274 ^ 1'h1;
  assign T274 = T275 | io_in_3_valid;
  assign T275 = T276 | io_in_2_valid;
  assign T276 = T277 | io_in_1_valid;
  assign T277 = T278 | io_in_0_valid;
  assign T278 = T279 | T192;
  assign T279 = T280 | T195;
  assign T280 = T281 | T198;
  assign T281 = T282 | T201;
  assign T282 = T283 | T204;
  assign T283 = T284 | T207;
  assign T284 = T212 | T210;
  assign T285 = T287 & T286;
  assign T286 = last_grant < 3'h4;
  assign T287 = T288 ^ 1'h1;
  assign T288 = T289 | T204;
  assign T289 = T290 | T207;
  assign T290 = T212 | T210;
  assign T291 = lockIdx == 3'h4;
  assign io_in_5_ready = T292;
  assign T292 = T293 & io_out_ready;
  assign T293 = locked ? T315 : T294;
  assign T294 = T308 | T295;
  assign T295 = T296 ^ 1'h1;
  assign T296 = T297 | io_in_4_valid;
  assign T297 = T298 | io_in_3_valid;
  assign T298 = T299 | io_in_2_valid;
  assign T299 = T300 | io_in_1_valid;
  assign T300 = T301 | io_in_0_valid;
  assign T301 = T302 | T192;
  assign T302 = T303 | T195;
  assign T303 = T304 | T198;
  assign T304 = T305 | T201;
  assign T305 = T306 | T204;
  assign T306 = T307 | T207;
  assign T307 = T212 | T210;
  assign T308 = T310 & T309;
  assign T309 = last_grant < 3'h5;
  assign T310 = T311 ^ 1'h1;
  assign T311 = T312 | T201;
  assign T312 = T313 | T204;
  assign T313 = T314 | T207;
  assign T314 = T212 | T210;
  assign T315 = lockIdx == 3'h5;
  assign io_in_6_ready = T316;
  assign T316 = T317 & io_out_ready;
  assign T317 = locked ? T341 : T318;
  assign T318 = T333 | T319;
  assign T319 = T320 ^ 1'h1;
  assign T320 = T321 | io_in_5_valid;
  assign T321 = T322 | io_in_4_valid;
  assign T322 = T323 | io_in_3_valid;
  assign T323 = T324 | io_in_2_valid;
  assign T324 = T325 | io_in_1_valid;
  assign T325 = T326 | io_in_0_valid;
  assign T326 = T327 | T192;
  assign T327 = T328 | T195;
  assign T328 = T329 | T198;
  assign T329 = T330 | T201;
  assign T330 = T331 | T204;
  assign T331 = T332 | T207;
  assign T332 = T212 | T210;
  assign T333 = T335 & T334;
  assign T334 = last_grant < 3'h6;
  assign T335 = T336 ^ 1'h1;
  assign T336 = T337 | T198;
  assign T337 = T338 | T201;
  assign T338 = T339 | T204;
  assign T339 = T340 | T207;
  assign T340 = T212 | T210;
  assign T341 = lockIdx == 3'h6;
  assign io_in_7_ready = T342;
  assign T342 = T343 & io_out_ready;
  assign T343 = locked ? T369 : T344;
  assign T344 = T360 | T345;
  assign T345 = T346 ^ 1'h1;
  assign T346 = T347 | io_in_6_valid;
  assign T347 = T348 | io_in_5_valid;
  assign T348 = T349 | io_in_4_valid;
  assign T349 = T350 | io_in_3_valid;
  assign T350 = T351 | io_in_2_valid;
  assign T351 = T352 | io_in_1_valid;
  assign T352 = T353 | io_in_0_valid;
  assign T353 = T354 | T192;
  assign T354 = T355 | T195;
  assign T355 = T356 | T198;
  assign T356 = T357 | T201;
  assign T357 = T358 | T204;
  assign T358 = T359 | T207;
  assign T359 = T212 | T210;
  assign T360 = T362 & T361;
  assign T361 = last_grant < 3'h7;
  assign T362 = T363 ^ 1'h1;
  assign T363 = T364 | T195;
  assign T364 = T365 | T198;
  assign T365 = T366 | T201;
  assign T366 = T367 | T204;
  assign T367 = T368 | T207;
  assign T368 = T212 | T210;
  assign T369 = lockIdx == 3'h7;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T17) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h7;
    end else if(T45) begin
      lockIdx <= T31;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T55) begin
      locked <= 1'h0;
    end else if(T45) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R58 <= 2'h0;
    end else if(T47) begin
      R58 <= T57;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input  io_in_7_bits_payload_manager_xact_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input  io_in_6_bits_payload_manager_xact_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input  io_in_5_bits_payload_manager_xact_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input  io_in_4_bits_payload_manager_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input  io_in_3_bits_payload_manager_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input  io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input  io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input  io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output io_out_bits_payload_manager_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  reg [2:0] last_grant;
  wire[2:0] T253;
  wire[2:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire T53;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T27 ? 3'h1 : T0;
  assign T0 = T25 ? 3'h2 : T1;
  assign T1 = T23 ? 3'h3 : T2;
  assign T2 = T21 ? 3'h4 : T3;
  assign T3 = T19 ? 3'h5 : T4;
  assign T4 = T17 ? 3'h6 : T5;
  assign T5 = T13 ? 3'h7 : T6;
  assign T6 = io_in_0_valid ? 3'h0 : T7;
  assign T7 = io_in_1_valid ? 3'h1 : T8;
  assign T8 = io_in_2_valid ? 3'h2 : T9;
  assign T9 = io_in_3_valid ? 3'h3 : T10;
  assign T10 = io_in_4_valid ? 3'h4 : T11;
  assign T11 = io_in_5_valid ? 3'h5 : T12;
  assign T12 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T13 = io_in_7_valid & T14;
  assign T14 = last_grant < 3'h7;
  assign T253 = reset ? 3'h0 : T15;
  assign T15 = T16 ? chosen : last_grant;
  assign T16 = io_out_ready & io_out_valid;
  assign T17 = io_in_6_valid & T18;
  assign T18 = last_grant < 3'h6;
  assign T19 = io_in_5_valid & T20;
  assign T20 = last_grant < 3'h5;
  assign T21 = io_in_4_valid & T22;
  assign T22 = last_grant < 3'h4;
  assign T23 = io_in_3_valid & T24;
  assign T24 = last_grant < 3'h3;
  assign T25 = io_in_2_valid & T26;
  assign T26 = last_grant < 3'h2;
  assign T27 = io_in_1_valid & T28;
  assign T28 = last_grant < 3'h1;
  assign io_out_bits_payload_manager_xact_id = T29;
  assign T29 = T43 ? T37 : T30;
  assign T30 = T36 ? T34 : T31;
  assign T31 = T32 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T32 = T33[1'h0:1'h0];
  assign T33 = chosen;
  assign T34 = T35 ? io_in_3_bits_payload_manager_xact_id : io_in_2_bits_payload_manager_xact_id;
  assign T35 = T33[1'h0:1'h0];
  assign T36 = T33[1'h1:1'h1];
  assign T37 = T42 ? T40 : T38;
  assign T38 = T39 ? io_in_5_bits_payload_manager_xact_id : io_in_4_bits_payload_manager_xact_id;
  assign T39 = T33[1'h0:1'h0];
  assign T40 = T41 ? io_in_7_bits_payload_manager_xact_id : io_in_6_bits_payload_manager_xact_id;
  assign T41 = T33[1'h0:1'h0];
  assign T42 = T33[1'h1:1'h1];
  assign T43 = T33[2'h2:2'h2];
  assign io_out_bits_header_dst = T44;
  assign T44 = T57 ? T51 : T45;
  assign T45 = T50 ? T48 : T46;
  assign T46 = T47 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T47 = T33[1'h0:1'h0];
  assign T48 = T49 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T49 = T33[1'h0:1'h0];
  assign T50 = T33[1'h1:1'h1];
  assign T51 = T56 ? T54 : T52;
  assign T52 = T53 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T53 = T33[1'h0:1'h0];
  assign T54 = T55 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T55 = T33[1'h0:1'h0];
  assign T56 = T33[1'h1:1'h1];
  assign T57 = T33[2'h2:2'h2];
  assign io_out_bits_header_src = T58;
  assign T58 = T71 ? T65 : T59;
  assign T59 = T64 ? T62 : T60;
  assign T60 = T61 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T61 = T33[1'h0:1'h0];
  assign T62 = T63 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T63 = T33[1'h0:1'h0];
  assign T64 = T33[1'h1:1'h1];
  assign T65 = T70 ? T68 : T66;
  assign T66 = T67 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T67 = T33[1'h0:1'h0];
  assign T68 = T69 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T69 = T33[1'h0:1'h0];
  assign T70 = T33[1'h1:1'h1];
  assign T71 = T33[2'h2:2'h2];
  assign io_out_valid = T72;
  assign T72 = T85 ? T79 : T73;
  assign T73 = T78 ? T76 : T74;
  assign T74 = T75 ? io_in_1_valid : io_in_0_valid;
  assign T75 = T33[1'h0:1'h0];
  assign T76 = T77 ? io_in_3_valid : io_in_2_valid;
  assign T77 = T33[1'h0:1'h0];
  assign T78 = T33[1'h1:1'h1];
  assign T79 = T84 ? T82 : T80;
  assign T80 = T81 ? io_in_5_valid : io_in_4_valid;
  assign T81 = T33[1'h0:1'h0];
  assign T82 = T83 ? io_in_7_valid : io_in_6_valid;
  assign T83 = T33[1'h0:1'h0];
  assign T84 = T33[1'h1:1'h1];
  assign T85 = T33[2'h2:2'h2];
  assign io_in_0_ready = T86;
  assign T86 = T87 & io_out_ready;
  assign T87 = T112 | T88;
  assign T88 = T89 ^ 1'h1;
  assign T89 = T92 | T90;
  assign T90 = io_in_7_valid & T91;
  assign T91 = last_grant < 3'h7;
  assign T92 = T95 | T93;
  assign T93 = io_in_6_valid & T94;
  assign T94 = last_grant < 3'h6;
  assign T95 = T98 | T96;
  assign T96 = io_in_5_valid & T97;
  assign T97 = last_grant < 3'h5;
  assign T98 = T101 | T99;
  assign T99 = io_in_4_valid & T100;
  assign T100 = last_grant < 3'h4;
  assign T101 = T104 | T102;
  assign T102 = io_in_3_valid & T103;
  assign T103 = last_grant < 3'h3;
  assign T104 = T107 | T105;
  assign T105 = io_in_2_valid & T106;
  assign T106 = last_grant < 3'h2;
  assign T107 = T110 | T108;
  assign T108 = io_in_1_valid & T109;
  assign T109 = last_grant < 3'h1;
  assign T110 = io_in_0_valid & T111;
  assign T111 = last_grant < 3'h0;
  assign T112 = last_grant < 3'h0;
  assign io_in_1_ready = T113;
  assign T113 = T114 & io_out_ready;
  assign T114 = T124 | T115;
  assign T115 = T116 ^ 1'h1;
  assign T116 = T117 | io_in_0_valid;
  assign T117 = T118 | T90;
  assign T118 = T119 | T93;
  assign T119 = T120 | T96;
  assign T120 = T121 | T99;
  assign T121 = T122 | T102;
  assign T122 = T123 | T105;
  assign T123 = T110 | T108;
  assign T124 = T126 & T125;
  assign T125 = last_grant < 3'h1;
  assign T126 = T110 ^ 1'h1;
  assign io_in_2_ready = T127;
  assign T127 = T128 & io_out_ready;
  assign T128 = T139 | T129;
  assign T129 = T130 ^ 1'h1;
  assign T130 = T131 | io_in_1_valid;
  assign T131 = T132 | io_in_0_valid;
  assign T132 = T133 | T90;
  assign T133 = T134 | T93;
  assign T134 = T135 | T96;
  assign T135 = T136 | T99;
  assign T136 = T137 | T102;
  assign T137 = T138 | T105;
  assign T138 = T110 | T108;
  assign T139 = T141 & T140;
  assign T140 = last_grant < 3'h2;
  assign T141 = T142 ^ 1'h1;
  assign T142 = T110 | T108;
  assign io_in_3_ready = T143;
  assign T143 = T144 & io_out_ready;
  assign T144 = T156 | T145;
  assign T145 = T146 ^ 1'h1;
  assign T146 = T147 | io_in_2_valid;
  assign T147 = T148 | io_in_1_valid;
  assign T148 = T149 | io_in_0_valid;
  assign T149 = T150 | T90;
  assign T150 = T151 | T93;
  assign T151 = T152 | T96;
  assign T152 = T153 | T99;
  assign T153 = T154 | T102;
  assign T154 = T155 | T105;
  assign T155 = T110 | T108;
  assign T156 = T158 & T157;
  assign T157 = last_grant < 3'h3;
  assign T158 = T159 ^ 1'h1;
  assign T159 = T160 | T105;
  assign T160 = T110 | T108;
  assign io_in_4_ready = T161;
  assign T161 = T162 & io_out_ready;
  assign T162 = T175 | T163;
  assign T163 = T164 ^ 1'h1;
  assign T164 = T165 | io_in_3_valid;
  assign T165 = T166 | io_in_2_valid;
  assign T166 = T167 | io_in_1_valid;
  assign T167 = T168 | io_in_0_valid;
  assign T168 = T169 | T90;
  assign T169 = T170 | T93;
  assign T170 = T171 | T96;
  assign T171 = T172 | T99;
  assign T172 = T173 | T102;
  assign T173 = T174 | T105;
  assign T174 = T110 | T108;
  assign T175 = T177 & T176;
  assign T176 = last_grant < 3'h4;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T179 | T102;
  assign T179 = T180 | T105;
  assign T180 = T110 | T108;
  assign io_in_5_ready = T181;
  assign T181 = T182 & io_out_ready;
  assign T182 = T196 | T183;
  assign T183 = T184 ^ 1'h1;
  assign T184 = T185 | io_in_4_valid;
  assign T185 = T186 | io_in_3_valid;
  assign T186 = T187 | io_in_2_valid;
  assign T187 = T188 | io_in_1_valid;
  assign T188 = T189 | io_in_0_valid;
  assign T189 = T190 | T90;
  assign T190 = T191 | T93;
  assign T191 = T192 | T96;
  assign T192 = T193 | T99;
  assign T193 = T194 | T102;
  assign T194 = T195 | T105;
  assign T195 = T110 | T108;
  assign T196 = T198 & T197;
  assign T197 = last_grant < 3'h5;
  assign T198 = T199 ^ 1'h1;
  assign T199 = T200 | T99;
  assign T200 = T201 | T102;
  assign T201 = T202 | T105;
  assign T202 = T110 | T108;
  assign io_in_6_ready = T203;
  assign T203 = T204 & io_out_ready;
  assign T204 = T219 | T205;
  assign T205 = T206 ^ 1'h1;
  assign T206 = T207 | io_in_5_valid;
  assign T207 = T208 | io_in_4_valid;
  assign T208 = T209 | io_in_3_valid;
  assign T209 = T210 | io_in_2_valid;
  assign T210 = T211 | io_in_1_valid;
  assign T211 = T212 | io_in_0_valid;
  assign T212 = T213 | T90;
  assign T213 = T214 | T93;
  assign T214 = T215 | T96;
  assign T215 = T216 | T99;
  assign T216 = T217 | T102;
  assign T217 = T218 | T105;
  assign T218 = T110 | T108;
  assign T219 = T221 & T220;
  assign T220 = last_grant < 3'h6;
  assign T221 = T222 ^ 1'h1;
  assign T222 = T223 | T96;
  assign T223 = T224 | T99;
  assign T224 = T225 | T102;
  assign T225 = T226 | T105;
  assign T226 = T110 | T108;
  assign io_in_7_ready = T227;
  assign T227 = T228 & io_out_ready;
  assign T228 = T244 | T229;
  assign T229 = T230 ^ 1'h1;
  assign T230 = T231 | io_in_6_valid;
  assign T231 = T232 | io_in_5_valid;
  assign T232 = T233 | io_in_4_valid;
  assign T233 = T234 | io_in_3_valid;
  assign T234 = T235 | io_in_2_valid;
  assign T235 = T236 | io_in_1_valid;
  assign T236 = T237 | io_in_0_valid;
  assign T237 = T238 | T90;
  assign T238 = T239 | T93;
  assign T239 = T240 | T96;
  assign T240 = T241 | T99;
  assign T241 = T242 | T102;
  assign T242 = T243 | T105;
  assign T243 = T110 | T108;
  assign T244 = T246 & T245;
  assign T245 = last_grant < 3'h7;
  assign T246 = T247 ^ 1'h1;
  assign T247 = T248 | T93;
  assign T248 = T249 | T96;
  assign T249 = T250 | T99;
  assign T250 = T251 | T102;
  assign T251 = T252 | T105;
  assign T252 = T110 | T108;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T16) begin
      last_grant <= chosen;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatPassesId(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [1:0] io_in_7_acquire_bits_header_src,
    input [1:0] io_in_7_acquire_bits_header_dst,
    input [25:0] io_in_7_acquire_bits_payload_addr,
    input [4:0] io_in_7_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_7_acquire_bits_payload_data,
    input  io_in_7_acquire_bits_payload_uncached,
    input [1:0] io_in_7_acquire_bits_payload_a_type,
    input [9:0] io_in_7_acquire_bits_payload_subblock,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_header_src,
    output[1:0] io_in_7_grant_bits_header_dst,
    output[3:0] io_in_7_grant_bits_payload_data,
    output[4:0] io_in_7_grant_bits_payload_client_xact_id,
    output io_in_7_grant_bits_payload_manager_xact_id,
    output io_in_7_grant_bits_payload_uncached,
    output[1:0] io_in_7_grant_bits_payload_g_type,
    output io_in_7_finish_ready,
    input  io_in_7_finish_valid,
    input [1:0] io_in_7_finish_bits_header_src,
    input [1:0] io_in_7_finish_bits_header_dst,
    input  io_in_7_finish_bits_payload_manager_xact_id,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [1:0] io_in_6_acquire_bits_header_src,
    input [1:0] io_in_6_acquire_bits_header_dst,
    input [25:0] io_in_6_acquire_bits_payload_addr,
    input [4:0] io_in_6_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_6_acquire_bits_payload_data,
    input  io_in_6_acquire_bits_payload_uncached,
    input [1:0] io_in_6_acquire_bits_payload_a_type,
    input [9:0] io_in_6_acquire_bits_payload_subblock,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_header_src,
    output[1:0] io_in_6_grant_bits_header_dst,
    output[3:0] io_in_6_grant_bits_payload_data,
    output[4:0] io_in_6_grant_bits_payload_client_xact_id,
    output io_in_6_grant_bits_payload_manager_xact_id,
    output io_in_6_grant_bits_payload_uncached,
    output[1:0] io_in_6_grant_bits_payload_g_type,
    output io_in_6_finish_ready,
    input  io_in_6_finish_valid,
    input [1:0] io_in_6_finish_bits_header_src,
    input [1:0] io_in_6_finish_bits_header_dst,
    input  io_in_6_finish_bits_payload_manager_xact_id,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [1:0] io_in_5_acquire_bits_header_src,
    input [1:0] io_in_5_acquire_bits_header_dst,
    input [25:0] io_in_5_acquire_bits_payload_addr,
    input [4:0] io_in_5_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_5_acquire_bits_payload_data,
    input  io_in_5_acquire_bits_payload_uncached,
    input [1:0] io_in_5_acquire_bits_payload_a_type,
    input [9:0] io_in_5_acquire_bits_payload_subblock,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_header_src,
    output[1:0] io_in_5_grant_bits_header_dst,
    output[3:0] io_in_5_grant_bits_payload_data,
    output[4:0] io_in_5_grant_bits_payload_client_xact_id,
    output io_in_5_grant_bits_payload_manager_xact_id,
    output io_in_5_grant_bits_payload_uncached,
    output[1:0] io_in_5_grant_bits_payload_g_type,
    output io_in_5_finish_ready,
    input  io_in_5_finish_valid,
    input [1:0] io_in_5_finish_bits_header_src,
    input [1:0] io_in_5_finish_bits_header_dst,
    input  io_in_5_finish_bits_payload_manager_xact_id,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [1:0] io_in_4_acquire_bits_header_src,
    input [1:0] io_in_4_acquire_bits_header_dst,
    input [25:0] io_in_4_acquire_bits_payload_addr,
    input [4:0] io_in_4_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_4_acquire_bits_payload_data,
    input  io_in_4_acquire_bits_payload_uncached,
    input [1:0] io_in_4_acquire_bits_payload_a_type,
    input [9:0] io_in_4_acquire_bits_payload_subblock,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_header_src,
    output[1:0] io_in_4_grant_bits_header_dst,
    output[3:0] io_in_4_grant_bits_payload_data,
    output[4:0] io_in_4_grant_bits_payload_client_xact_id,
    output io_in_4_grant_bits_payload_manager_xact_id,
    output io_in_4_grant_bits_payload_uncached,
    output[1:0] io_in_4_grant_bits_payload_g_type,
    output io_in_4_finish_ready,
    input  io_in_4_finish_valid,
    input [1:0] io_in_4_finish_bits_header_src,
    input [1:0] io_in_4_finish_bits_header_dst,
    input  io_in_4_finish_bits_payload_manager_xact_id,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [1:0] io_in_3_acquire_bits_header_src,
    input [1:0] io_in_3_acquire_bits_header_dst,
    input [25:0] io_in_3_acquire_bits_payload_addr,
    input [4:0] io_in_3_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_3_acquire_bits_payload_data,
    input  io_in_3_acquire_bits_payload_uncached,
    input [1:0] io_in_3_acquire_bits_payload_a_type,
    input [9:0] io_in_3_acquire_bits_payload_subblock,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_header_src,
    output[1:0] io_in_3_grant_bits_header_dst,
    output[3:0] io_in_3_grant_bits_payload_data,
    output[4:0] io_in_3_grant_bits_payload_client_xact_id,
    output io_in_3_grant_bits_payload_manager_xact_id,
    output io_in_3_grant_bits_payload_uncached,
    output[1:0] io_in_3_grant_bits_payload_g_type,
    output io_in_3_finish_ready,
    input  io_in_3_finish_valid,
    input [1:0] io_in_3_finish_bits_header_src,
    input [1:0] io_in_3_finish_bits_header_dst,
    input  io_in_3_finish_bits_payload_manager_xact_id,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [4:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_2_acquire_bits_payload_data,
    input  io_in_2_acquire_bits_payload_uncached,
    input [1:0] io_in_2_acquire_bits_payload_a_type,
    input [9:0] io_in_2_acquire_bits_payload_subblock,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[3:0] io_in_2_grant_bits_payload_data,
    output[4:0] io_in_2_grant_bits_payload_client_xact_id,
    output io_in_2_grant_bits_payload_manager_xact_id,
    output io_in_2_grant_bits_payload_uncached,
    output[1:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input  io_in_2_finish_bits_payload_manager_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [4:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_1_acquire_bits_payload_data,
    input  io_in_1_acquire_bits_payload_uncached,
    input [1:0] io_in_1_acquire_bits_payload_a_type,
    input [9:0] io_in_1_acquire_bits_payload_subblock,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[3:0] io_in_1_grant_bits_payload_data,
    output[4:0] io_in_1_grant_bits_payload_client_xact_id,
    output io_in_1_grant_bits_payload_manager_xact_id,
    output io_in_1_grant_bits_payload_uncached,
    output[1:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input  io_in_1_finish_bits_payload_manager_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [4:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [3:0] io_in_0_acquire_bits_payload_data,
    input  io_in_0_acquire_bits_payload_uncached,
    input [1:0] io_in_0_acquire_bits_payload_a_type,
    input [9:0] io_in_0_acquire_bits_payload_subblock,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[3:0] io_in_0_grant_bits_payload_data,
    output[4:0] io_in_0_grant_bits_payload_client_xact_id,
    output io_in_0_grant_bits_payload_manager_xact_id,
    output io_in_0_grant_bits_payload_uncached,
    output[1:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input  io_in_0_finish_bits_payload_manager_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[4:0] io_out_acquire_bits_payload_client_xact_id,
    output[3:0] io_out_acquire_bits_payload_data,
    output io_out_acquire_bits_payload_uncached,
    output[1:0] io_out_acquire_bits_payload_a_type,
    output[9:0] io_out_acquire_bits_payload_subblock,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [3:0] io_out_grant_bits_payload_data,
    input [4:0] io_out_grant_bits_payload_client_xact_id,
    input  io_out_grant_bits_payload_manager_xact_id,
    input  io_out_grant_bits_payload_uncached,
    input [1:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output io_out_finish_bits_payload_manager_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire LockingRRArbiter_24_io_in_7_ready;
  wire LockingRRArbiter_24_io_in_6_ready;
  wire LockingRRArbiter_24_io_in_5_ready;
  wire LockingRRArbiter_24_io_in_4_ready;
  wire LockingRRArbiter_24_io_in_3_ready;
  wire LockingRRArbiter_24_io_in_2_ready;
  wire LockingRRArbiter_24_io_in_1_ready;
  wire LockingRRArbiter_24_io_in_0_ready;
  wire LockingRRArbiter_24_io_out_valid;
  wire[1:0] LockingRRArbiter_24_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_24_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_24_io_out_bits_payload_addr;
  wire[4:0] LockingRRArbiter_24_io_out_bits_payload_client_xact_id;
  wire[3:0] LockingRRArbiter_24_io_out_bits_payload_data;
  wire LockingRRArbiter_24_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_24_io_out_bits_payload_a_type;
  wire[9:0] LockingRRArbiter_24_io_out_bits_payload_subblock;
  wire finish_arb_io_in_7_ready;
  wire finish_arb_io_in_6_ready;
  wire finish_arb_io_in_5_ready;
  wire finish_arb_io_in_4_ready;
  wire finish_arb_io_in_3_ready;
  wire finish_arb_io_in_2_ready;
  wire finish_arb_io_in_1_ready;
  wire finish_arb_io_in_0_ready;
  wire finish_arb_io_out_valid;
  wire[1:0] finish_arb_io_out_bits_header_src;
  wire[1:0] finish_arb_io_out_bits_header_dst;
  wire finish_arb_io_out_bits_payload_manager_xact_id;


  assign io_out_finish_bits_payload_manager_xact_id = finish_arb_io_out_bits_payload_manager_xact_id;
  assign io_out_finish_bits_header_dst = finish_arb_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = finish_arb_io_out_bits_header_src;
  assign io_out_finish_valid = finish_arb_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T15 ? io_in_7_grant_ready : T1;
  assign T1 = T14 ? io_in_6_grant_ready : T2;
  assign T2 = T13 ? io_in_5_grant_ready : T3;
  assign T3 = T12 ? io_in_4_grant_ready : T4;
  assign T4 = T11 ? io_in_3_grant_ready : T5;
  assign T5 = T10 ? io_in_2_grant_ready : T6;
  assign T6 = T9 ? io_in_1_grant_ready : T7;
  assign T7 = T8 ? io_in_0_grant_ready : 1'h0;
  assign T8 = io_out_grant_bits_payload_client_xact_id == 5'h0;
  assign T9 = io_out_grant_bits_payload_client_xact_id == 5'h1;
  assign T10 = io_out_grant_bits_payload_client_xact_id == 5'h2;
  assign T11 = io_out_grant_bits_payload_client_xact_id == 5'h3;
  assign T12 = io_out_grant_bits_payload_client_xact_id == 5'h4;
  assign T13 = io_out_grant_bits_payload_client_xact_id == 5'h5;
  assign T14 = io_out_grant_bits_payload_client_xact_id == 5'h6;
  assign T15 = io_out_grant_bits_payload_client_xact_id == 5'h7;
  assign io_out_acquire_bits_payload_subblock = LockingRRArbiter_24_io_out_bits_payload_subblock;
  assign io_out_acquire_bits_payload_a_type = LockingRRArbiter_24_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_uncached = LockingRRArbiter_24_io_out_bits_payload_uncached;
  assign io_out_acquire_bits_payload_data = LockingRRArbiter_24_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = LockingRRArbiter_24_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = LockingRRArbiter_24_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = LockingRRArbiter_24_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = LockingRRArbiter_24_io_out_bits_header_src;
  assign io_out_acquire_valid = LockingRRArbiter_24_io_out_valid;
  assign io_in_0_finish_ready = finish_arb_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_0_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T16;
  assign T16 = T8 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_24_io_in_0_ready;
  assign io_in_1_finish_ready = finish_arb_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_1_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_24_io_in_1_ready;
  assign io_in_2_finish_ready = finish_arb_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_2_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T18;
  assign T18 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = LockingRRArbiter_24_io_in_2_ready;
  assign io_in_3_finish_ready = finish_arb_io_in_3_ready;
  assign io_in_3_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_3_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_3_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_3_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_3_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_3_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_3_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_3_grant_valid = T19;
  assign T19 = T11 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = LockingRRArbiter_24_io_in_3_ready;
  assign io_in_4_finish_ready = finish_arb_io_in_4_ready;
  assign io_in_4_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_4_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_4_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_4_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_4_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_4_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_4_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_4_grant_valid = T20;
  assign T20 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = LockingRRArbiter_24_io_in_4_ready;
  assign io_in_5_finish_ready = finish_arb_io_in_5_ready;
  assign io_in_5_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_5_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_5_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_5_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_5_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_5_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_5_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_5_grant_valid = T21;
  assign T21 = T13 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = LockingRRArbiter_24_io_in_5_ready;
  assign io_in_6_finish_ready = finish_arb_io_in_6_ready;
  assign io_in_6_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_6_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_6_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_6_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_6_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_6_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_6_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_6_grant_valid = T22;
  assign T22 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = LockingRRArbiter_24_io_in_6_ready;
  assign io_in_7_finish_ready = finish_arb_io_in_7_ready;
  assign io_in_7_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_7_grant_bits_payload_uncached = io_out_grant_bits_payload_uncached;
  assign io_in_7_grant_bits_payload_manager_xact_id = io_out_grant_bits_payload_manager_xact_id;
  assign io_in_7_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_7_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_7_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_7_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_7_grant_valid = T23;
  assign T23 = T15 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = LockingRRArbiter_24_io_in_7_ready;
  LockingRRArbiter_14 LockingRRArbiter_24(.clk(clk), .reset(reset),
       .io_in_7_ready( LockingRRArbiter_24_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_header_src( io_in_7_acquire_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_acquire_bits_header_dst ),
       .io_in_7_bits_payload_addr( io_in_7_acquire_bits_payload_addr ),
       .io_in_7_bits_payload_client_xact_id( io_in_7_acquire_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_data( io_in_7_acquire_bits_payload_data ),
       .io_in_7_bits_payload_uncached( io_in_7_acquire_bits_payload_uncached ),
       .io_in_7_bits_payload_a_type( io_in_7_acquire_bits_payload_a_type ),
       .io_in_7_bits_payload_subblock( io_in_7_acquire_bits_payload_subblock ),
       .io_in_6_ready( LockingRRArbiter_24_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_header_src( io_in_6_acquire_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_acquire_bits_header_dst ),
       .io_in_6_bits_payload_addr( io_in_6_acquire_bits_payload_addr ),
       .io_in_6_bits_payload_client_xact_id( io_in_6_acquire_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_data( io_in_6_acquire_bits_payload_data ),
       .io_in_6_bits_payload_uncached( io_in_6_acquire_bits_payload_uncached ),
       .io_in_6_bits_payload_a_type( io_in_6_acquire_bits_payload_a_type ),
       .io_in_6_bits_payload_subblock( io_in_6_acquire_bits_payload_subblock ),
       .io_in_5_ready( LockingRRArbiter_24_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_header_src( io_in_5_acquire_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_acquire_bits_header_dst ),
       .io_in_5_bits_payload_addr( io_in_5_acquire_bits_payload_addr ),
       .io_in_5_bits_payload_client_xact_id( io_in_5_acquire_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_data( io_in_5_acquire_bits_payload_data ),
       .io_in_5_bits_payload_uncached( io_in_5_acquire_bits_payload_uncached ),
       .io_in_5_bits_payload_a_type( io_in_5_acquire_bits_payload_a_type ),
       .io_in_5_bits_payload_subblock( io_in_5_acquire_bits_payload_subblock ),
       .io_in_4_ready( LockingRRArbiter_24_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_header_src( io_in_4_acquire_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_acquire_bits_header_dst ),
       .io_in_4_bits_payload_addr( io_in_4_acquire_bits_payload_addr ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_acquire_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_data( io_in_4_acquire_bits_payload_data ),
       .io_in_4_bits_payload_uncached( io_in_4_acquire_bits_payload_uncached ),
       .io_in_4_bits_payload_a_type( io_in_4_acquire_bits_payload_a_type ),
       .io_in_4_bits_payload_subblock( io_in_4_acquire_bits_payload_subblock ),
       .io_in_3_ready( LockingRRArbiter_24_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_header_src( io_in_3_acquire_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_acquire_bits_header_dst ),
       .io_in_3_bits_payload_addr( io_in_3_acquire_bits_payload_addr ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_acquire_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_data( io_in_3_acquire_bits_payload_data ),
       .io_in_3_bits_payload_uncached( io_in_3_acquire_bits_payload_uncached ),
       .io_in_3_bits_payload_a_type( io_in_3_acquire_bits_payload_a_type ),
       .io_in_3_bits_payload_subblock( io_in_3_acquire_bits_payload_subblock ),
       .io_in_2_ready( LockingRRArbiter_24_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_uncached( io_in_2_acquire_bits_payload_uncached ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_subblock( io_in_2_acquire_bits_payload_subblock ),
       .io_in_1_ready( LockingRRArbiter_24_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_uncached( io_in_1_acquire_bits_payload_uncached ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_subblock( io_in_1_acquire_bits_payload_subblock ),
       .io_in_0_ready( LockingRRArbiter_24_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_uncached( io_in_0_acquire_bits_payload_uncached ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_subblock( io_in_0_acquire_bits_payload_subblock ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_24_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_24_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_24_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_24_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_24_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_24_io_out_bits_payload_data ),
       .io_out_bits_payload_uncached( LockingRRArbiter_24_io_out_bits_payload_uncached ),
       .io_out_bits_payload_a_type( LockingRRArbiter_24_io_out_bits_payload_a_type ),
       .io_out_bits_payload_subblock( LockingRRArbiter_24_io_out_bits_payload_subblock )
       //.io_chosen(  )
  );
  RRArbiter_2 finish_arb(.clk(clk), .reset(reset),
       .io_in_7_ready( finish_arb_io_in_7_ready ),
       .io_in_7_valid( io_in_7_finish_valid ),
       .io_in_7_bits_header_src( io_in_7_finish_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_finish_bits_header_dst ),
       .io_in_7_bits_payload_manager_xact_id( io_in_7_finish_bits_payload_manager_xact_id ),
       .io_in_6_ready( finish_arb_io_in_6_ready ),
       .io_in_6_valid( io_in_6_finish_valid ),
       .io_in_6_bits_header_src( io_in_6_finish_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_finish_bits_header_dst ),
       .io_in_6_bits_payload_manager_xact_id( io_in_6_finish_bits_payload_manager_xact_id ),
       .io_in_5_ready( finish_arb_io_in_5_ready ),
       .io_in_5_valid( io_in_5_finish_valid ),
       .io_in_5_bits_header_src( io_in_5_finish_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_finish_bits_header_dst ),
       .io_in_5_bits_payload_manager_xact_id( io_in_5_finish_bits_payload_manager_xact_id ),
       .io_in_4_ready( finish_arb_io_in_4_ready ),
       .io_in_4_valid( io_in_4_finish_valid ),
       .io_in_4_bits_header_src( io_in_4_finish_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_finish_bits_header_dst ),
       .io_in_4_bits_payload_manager_xact_id( io_in_4_finish_bits_payload_manager_xact_id ),
       .io_in_3_ready( finish_arb_io_in_3_ready ),
       .io_in_3_valid( io_in_3_finish_valid ),
       .io_in_3_bits_header_src( io_in_3_finish_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_finish_bits_header_dst ),
       .io_in_3_bits_payload_manager_xact_id( io_in_3_finish_bits_payload_manager_xact_id ),
       .io_in_2_ready( finish_arb_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( io_in_2_finish_bits_payload_manager_xact_id ),
       .io_in_1_ready( finish_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( io_in_1_finish_bits_payload_manager_xact_id ),
       .io_in_0_ready( finish_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( io_in_0_finish_bits_payload_manager_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( finish_arb_io_out_valid ),
       .io_out_bits_header_src( finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( finish_arb_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module L2BroadcastHub(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [135:0] io_inner_acquire_bits_payload_data,
    input  io_inner_acquire_bits_payload_uncached,
    input [1:0] io_inner_acquire_bits_payload_a_type,
    input [128:0] io_inner_acquire_bits_payload_subblock,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[135:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_manager_xact_id,
    output io_inner_grant_bits_payload_uncached,
    output[1:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [135:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    output[1:0] io_outer_acquire_bits_header_dst,
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[4:0] io_outer_acquire_bits_payload_client_xact_id,
    output[135:0] io_outer_acquire_bits_payload_data,
    output io_outer_acquire_bits_payload_uncached,
    output[1:0] io_outer_acquire_bits_payload_a_type,
    output[128:0] io_outer_acquire_bits_payload_subblock,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [135:0] io_outer_grant_bits_payload_data,
    input [4:0] io_outer_grant_bits_payload_client_xact_id,
    input  io_outer_grant_bits_payload_manager_xact_id,
    input  io_outer_grant_bits_payload_uncached,
    input [1:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    output io_outer_finish_valid,
    output[1:0] io_outer_finish_bits_header_src,
    output[1:0] io_outer_finish_bits_header_dst,
    output io_outer_finish_bits_payload_manager_xact_id,
    input  io_incoherent_1,
    input  io_incoherent_0
);

  wire[3:0] T222;
  wire[135:0] T223;
  wire[135:0] T224;
  wire[135:0] T225;
  wire[135:0] T226;
  wire[135:0] T227;
  wire[135:0] T228;
  wire[135:0] T229;
  wire[135:0] T230;
  wire T0;
  wire T1;
  wire any_acquire_conflict;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire sdq_rdy;
  wire T9;
  reg [3:0] sdq_val;
  wire[3:0] T231;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T232;
  wire sdq_enq;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[3:0] T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire[3:0] T233;
  wire free_sdq;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[3:0] T41;
  wire[1:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire[2:0] release_idx;
  wire[2:0] T52;
  wire[2:0] T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire[2:0] T57;
  wire[9:0] T234;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire T238;
  wire[3:0] T62;
  wire T239;
  wire T240;
  wire[1:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire[9:0] T241;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire[3:0] T75;
  wire[3:0] T76;
  wire[1:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire[9:0] T242;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[3:0] T86;
  wire[3:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire[9:0] T243;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire[1:0] T99;
  wire[1:0] T100;
  wire T101;
  wire T102;
  wire[9:0] T244;
  wire[3:0] T103;
  wire[3:0] T104;
  wire[1:0] T105;
  wire[1:0] T106;
  wire[1:0] T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire[9:0] T245;
  wire[3:0] T114;
  wire[3:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[3:0] T119;
  wire[3:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire T124;
  wire[9:0] T246;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[1:0] T127;
  wire[1:0] T128;
  wire[1:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  reg [1:0] rel_data_cnt;
  wire[1:0] T247;
  wire[1:0] T134;
  wire[1:0] T135;
  wire vwbdq_enq;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire voluntary;
  wire T144;
  wire T145;
  wire T146;
  wire[9:0] T248;
  wire[3:0] T147;
  wire[3:0] T148;
  wire[1:0] T149;
  wire[1:0] T150;
  wire[128:0] T249;
  wire[135:0] T151;
  wire[135:0] T152;
  wire[135:0] T153;
  wire[135:0] T154;
  reg [135:0] vwbdq_0;
  wire[135:0] T155;
  wire T156;
  wire T157;
  wire[3:0] T158;
  wire[1:0] T159;
  reg [135:0] vwbdq_1;
  wire[135:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire[1:0] T164;
  wire[135:0] T165;
  reg [135:0] vwbdq_2;
  wire[135:0] T166;
  wire T167;
  wire T168;
  reg [135:0] vwbdq_3;
  wire[135:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[135:0] T175;
  wire[135:0] T176;
  reg [135:0] sdq_0;
  wire[135:0] T177;
  wire T178;
  wire T179;
  wire[3:0] T180;
  wire[1:0] T181;
  reg [135:0] sdq_1;
  wire[135:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire[1:0] T186;
  wire[135:0] T187;
  reg [135:0] sdq_2;
  wire[135:0] T188;
  wire T189;
  wire T190;
  reg [135:0] sdq_3;
  wire[135:0] T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire[2:0] T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire VoluntaryReleaseTracker_io_inner_acquire_ready;
  wire VoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_src;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_dst;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_data;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_manager_xact_id;
  wire VoluntaryReleaseTracker_io_inner_grant_bits_payload_uncached;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type;
  wire VoluntaryReleaseTracker_io_inner_probe_valid;
  wire VoluntaryReleaseTracker_io_inner_release_ready;
  wire VoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[25:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr;
  wire[4:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data;
  wire VoluntaryReleaseTracker_io_outer_acquire_bits_payload_uncached;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type;
  wire[9:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subblock;
  wire VoluntaryReleaseTracker_io_outer_grant_ready;
  wire VoluntaryReleaseTracker_io_has_acquire_conflict;
  wire VoluntaryReleaseTracker_io_has_release_match;
  wire AcquireTracker_0_io_inner_acquire_ready;
  wire AcquireTracker_0_io_inner_grant_valid;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_0_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_0_io_inner_probe_valid;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_0_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_0_io_inner_release_ready;
  wire AcquireTracker_0_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_0_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_0_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_0_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_0_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_0_io_outer_grant_ready;
  wire AcquireTracker_0_io_has_acquire_conflict;
  wire AcquireTracker_0_io_has_release_match;
  wire AcquireTracker_1_io_inner_acquire_ready;
  wire AcquireTracker_1_io_inner_grant_valid;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_1_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_1_io_inner_probe_valid;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_1_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_1_io_inner_release_ready;
  wire AcquireTracker_1_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_1_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_1_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_1_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_1_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_1_io_outer_grant_ready;
  wire AcquireTracker_1_io_has_acquire_conflict;
  wire AcquireTracker_1_io_has_release_match;
  wire AcquireTracker_2_io_inner_acquire_ready;
  wire AcquireTracker_2_io_inner_grant_valid;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_2_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_2_io_inner_probe_valid;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_2_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_2_io_inner_release_ready;
  wire AcquireTracker_2_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_2_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_2_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_2_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_2_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_2_io_outer_grant_ready;
  wire AcquireTracker_2_io_has_acquire_conflict;
  wire AcquireTracker_2_io_has_release_match;
  wire AcquireTracker_3_io_inner_acquire_ready;
  wire AcquireTracker_3_io_inner_grant_valid;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_3_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_3_io_inner_probe_valid;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_3_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_3_io_inner_release_ready;
  wire AcquireTracker_3_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_3_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_3_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_3_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_3_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_3_io_outer_grant_ready;
  wire AcquireTracker_3_io_has_acquire_conflict;
  wire AcquireTracker_3_io_has_release_match;
  wire AcquireTracker_4_io_inner_acquire_ready;
  wire AcquireTracker_4_io_inner_grant_valid;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_4_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_4_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_4_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_4_io_inner_probe_valid;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_4_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_4_io_inner_release_ready;
  wire AcquireTracker_4_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_4_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_4_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_4_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_4_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_4_io_outer_grant_ready;
  wire AcquireTracker_4_io_has_acquire_conflict;
  wire AcquireTracker_4_io_has_release_match;
  wire AcquireTracker_5_io_inner_acquire_ready;
  wire AcquireTracker_5_io_inner_grant_valid;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_5_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_5_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_5_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_5_io_inner_probe_valid;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_5_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_5_io_inner_release_ready;
  wire AcquireTracker_5_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_5_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_5_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_5_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_5_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_5_io_outer_grant_ready;
  wire AcquireTracker_5_io_has_acquire_conflict;
  wire AcquireTracker_5_io_has_release_match;
  wire AcquireTracker_6_io_inner_acquire_ready;
  wire AcquireTracker_6_io_inner_grant_valid;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_dst;
  wire[3:0] AcquireTracker_6_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_6_io_inner_grant_bits_payload_manager_xact_id;
  wire AcquireTracker_6_io_inner_grant_bits_payload_uncached;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_6_io_inner_probe_valid;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_6_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_6_io_inner_release_ready;
  wire AcquireTracker_6_io_outer_acquire_valid;
  wire[25:0] AcquireTracker_6_io_outer_acquire_bits_payload_addr;
  wire[4:0] AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id;
  wire[3:0] AcquireTracker_6_io_outer_acquire_bits_payload_data;
  wire AcquireTracker_6_io_outer_acquire_bits_payload_uncached;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_payload_a_type;
  wire[9:0] AcquireTracker_6_io_outer_acquire_bits_payload_subblock;
  wire AcquireTracker_6_io_outer_grant_ready;
  wire AcquireTracker_6_io_has_acquire_conflict;
  wire alloc_arb_io_in_7_ready;
  wire alloc_arb_io_in_6_ready;
  wire alloc_arb_io_in_5_ready;
  wire alloc_arb_io_in_4_ready;
  wire alloc_arb_io_in_3_ready;
  wire alloc_arb_io_in_2_ready;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire probe_arb_io_in_7_ready;
  wire probe_arb_io_in_6_ready;
  wire probe_arb_io_in_5_ready;
  wire probe_arb_io_in_4_ready;
  wire probe_arb_io_in_3_ready;
  wire probe_arb_io_in_2_ready;
  wire probe_arb_io_in_1_ready;
  wire probe_arb_io_in_0_ready;
  wire probe_arb_io_out_valid;
  wire[1:0] probe_arb_io_out_bits_header_src;
  wire[1:0] probe_arb_io_out_bits_header_dst;
  wire[25:0] probe_arb_io_out_bits_payload_addr;
  wire[1:0] probe_arb_io_out_bits_payload_p_type;
  wire grant_arb_io_in_7_ready;
  wire grant_arb_io_in_6_ready;
  wire grant_arb_io_in_5_ready;
  wire grant_arb_io_in_4_ready;
  wire grant_arb_io_in_3_ready;
  wire grant_arb_io_in_2_ready;
  wire grant_arb_io_in_1_ready;
  wire grant_arb_io_in_0_ready;
  wire grant_arb_io_out_valid;
  wire[1:0] grant_arb_io_out_bits_header_src;
  wire[1:0] grant_arb_io_out_bits_header_dst;
  wire[1:0] grant_arb_io_out_bits_payload_client_xact_id;
  wire[3:0] grant_arb_io_out_bits_payload_manager_xact_id;
  wire grant_arb_io_out_bits_payload_uncached;
  wire[1:0] grant_arb_io_out_bits_payload_g_type;
  wire outer_arb_io_in_7_acquire_ready;
  wire outer_arb_io_in_7_grant_valid;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_7_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_7_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_7_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_7_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_7_grant_bits_payload_g_type;
  wire outer_arb_io_in_7_finish_ready;
  wire outer_arb_io_in_6_acquire_ready;
  wire outer_arb_io_in_6_grant_valid;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_6_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_6_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_6_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_6_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_6_grant_bits_payload_g_type;
  wire outer_arb_io_in_6_finish_ready;
  wire outer_arb_io_in_5_acquire_ready;
  wire outer_arb_io_in_5_grant_valid;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_5_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_5_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_5_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_5_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_5_grant_bits_payload_g_type;
  wire outer_arb_io_in_5_finish_ready;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_4_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_4_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_4_grant_bits_payload_g_type;
  wire outer_arb_io_in_4_finish_ready;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_3_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_3_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_3_grant_bits_payload_g_type;
  wire outer_arb_io_in_3_finish_ready;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_2_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_2_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_2_grant_bits_payload_g_type;
  wire outer_arb_io_in_2_finish_ready;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_1_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_1_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_1_grant_bits_payload_g_type;
  wire outer_arb_io_in_1_finish_ready;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_dst;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_data;
  wire[4:0] outer_arb_io_in_0_grant_bits_payload_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_payload_manager_xact_id;
  wire outer_arb_io_in_0_grant_bits_payload_uncached;
  wire[1:0] outer_arb_io_in_0_grant_bits_payload_g_type;
  wire outer_arb_io_in_0_finish_ready;
  wire outer_arb_io_out_acquire_valid;
  wire[1:0] outer_arb_io_out_acquire_bits_header_src;
  wire[1:0] outer_arb_io_out_acquire_bits_header_dst;
  wire[25:0] outer_arb_io_out_acquire_bits_payload_addr;
  wire[4:0] outer_arb_io_out_acquire_bits_payload_client_xact_id;
  wire[3:0] outer_arb_io_out_acquire_bits_payload_data;
  wire outer_arb_io_out_acquire_bits_payload_uncached;
  wire[1:0] outer_arb_io_out_acquire_bits_payload_a_type;
  wire[9:0] outer_arb_io_out_acquire_bits_payload_subblock;
  wire outer_arb_io_out_grant_ready;
  wire outer_arb_io_out_finish_valid;
  wire[1:0] outer_arb_io_out_finish_bits_header_src;
  wire[1:0] outer_arb_io_out_finish_bits_header_dst;
  wire outer_arb_io_out_finish_bits_payload_manager_xact_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    rel_data_cnt = {1{$random}};
    vwbdq_0 = {5{$random}};
    vwbdq_1 = {5{$random}};
    vwbdq_2 = {5{$random}};
    vwbdq_3 = {5{$random}};
    sdq_0 = {5{$random}};
    sdq_1 = {5{$random}};
    sdq_2 = {5{$random}};
    sdq_3 = {5{$random}};
  end
// synthesis translate_on
`endif

  assign T222 = io_outer_grant_bits_payload_data[2'h3:1'h0];
  assign T223 = {132'h0, VoluntaryReleaseTracker_io_inner_grant_bits_payload_data};
  assign T224 = {132'h0, AcquireTracker_0_io_inner_grant_bits_payload_data};
  assign T225 = {132'h0, AcquireTracker_1_io_inner_grant_bits_payload_data};
  assign T226 = {132'h0, AcquireTracker_2_io_inner_grant_bits_payload_data};
  assign T227 = {132'h0, AcquireTracker_3_io_inner_grant_bits_payload_data};
  assign T228 = {132'h0, AcquireTracker_4_io_inner_grant_bits_payload_data};
  assign T229 = {132'h0, AcquireTracker_5_io_inner_grant_bits_payload_data};
  assign T230 = {132'h0, AcquireTracker_6_io_inner_grant_bits_payload_data};
  assign T0 = T8 & T1;
  assign T1 = any_acquire_conflict ^ 1'h1;
  assign any_acquire_conflict = T2 | AcquireTracker_6_io_has_acquire_conflict;
  assign T2 = T3 | AcquireTracker_5_io_has_acquire_conflict;
  assign T3 = T4 | AcquireTracker_4_io_has_acquire_conflict;
  assign T4 = T5 | AcquireTracker_3_io_has_acquire_conflict;
  assign T5 = T6 | AcquireTracker_2_io_has_acquire_conflict;
  assign T6 = T7 | AcquireTracker_1_io_has_acquire_conflict;
  assign T7 = VoluntaryReleaseTracker_io_has_acquire_conflict | AcquireTracker_0_io_has_acquire_conflict;
  assign T8 = io_inner_acquire_valid & sdq_rdy;
  assign sdq_rdy = T9 ^ 1'h1;
  assign T9 = sdq_val == 4'hf;
  assign T231 = reset ? 4'h0 : T10;
  assign T10 = T43 ? T11 : sdq_val;
  assign T11 = T29 | T12;
  assign T12 = T19 & T13;
  assign T13 = 4'h0 - T232;
  assign T232 = {3'h0, sdq_enq};
  assign sdq_enq = T18 & T14;
  assign T14 = io_inner_acquire_bits_payload_uncached ? T15 : 1'h0;
  assign T15 = T17 | T16;
  assign T16 = 2'h2 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 2'h1 == io_inner_acquire_bits_payload_a_type;
  assign T18 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T19 = T28 ? 4'h1 : T20;
  assign T20 = T27 ? 4'h2 : T21;
  assign T21 = T26 ? 4'h4 : T22;
  assign T22 = T23 ? 4'h8 : 4'h0;
  assign T23 = T24[2'h3:2'h3];
  assign T24 = ~ T25;
  assign T25 = sdq_val[2'h3:1'h0];
  assign T26 = T24[2'h2:2'h2];
  assign T27 = T24[1'h1:1'h1];
  assign T28 = T24[1'h0:1'h0];
  assign T29 = sdq_val & T30;
  assign T30 = ~ T31;
  assign T31 = T41 & T32;
  assign T32 = 4'h0 - T233;
  assign T233 = {3'h0, free_sdq};
  assign free_sdq = T35 & T33;
  assign T33 = T34 == 2'h0;
  assign T34 = outer_arb_io_out_acquire_bits_payload_data[1'h1:1'h0];
  assign T35 = T40 & T36;
  assign T36 = io_outer_acquire_bits_payload_uncached ? T37 : 1'h0;
  assign T37 = T39 | T38;
  assign T38 = 2'h2 == io_outer_acquire_bits_payload_a_type;
  assign T39 = 2'h1 == io_outer_acquire_bits_payload_a_type;
  assign T40 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T41 = 1'h1 << T42;
  assign T42 = outer_arb_io_out_acquire_bits_payload_data[2'h3:2'h2];
  assign T43 = io_outer_acquire_valid | sdq_enq;
  assign T44 = T45;
  assign T45 = {io_incoherent_1, io_incoherent_0};
  assign T46 = T47;
  assign T47 = {T49, T48};
  assign T48 = 2'h2;
  assign T49 = 2'h0;
  assign T50 = io_inner_release_valid & T51;
  assign T51 = release_idx == 3'h7;
  assign release_idx = VoluntaryReleaseTracker_io_has_release_match ? 3'h0 : T52;
  assign T52 = AcquireTracker_0_io_has_release_match ? 3'h1 : T53;
  assign T53 = AcquireTracker_1_io_has_release_match ? 3'h2 : T54;
  assign T54 = AcquireTracker_2_io_has_release_match ? 3'h3 : T55;
  assign T55 = AcquireTracker_3_io_has_release_match ? 3'h4 : T56;
  assign T56 = AcquireTracker_4_io_has_release_match ? 3'h5 : T57;
  assign T57 = AcquireTracker_5_io_has_release_match ? 3'h6 : 3'h7;
  assign T234 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T58 = T59;
  assign T59 = {T61, T60};
  assign T60 = 2'h0;
  assign T61 = T235;
  assign T235 = T240 ? 1'h0 : T236;
  assign T236 = T239 ? 1'h1 : T237;
  assign T237 = T238 ? 2'h2 : 2'h3;
  assign T238 = T62[2'h2:2'h2];
  assign T62 = ~ sdq_val;
  assign T239 = T62[1'h1:1'h1];
  assign T240 = T62[1'h0:1'h0];
  assign T63 = T45;
  assign T64 = T65;
  assign T65 = {T67, T66};
  assign T66 = 2'h2;
  assign T67 = 2'h0;
  assign T68 = io_inner_release_valid & T69;
  assign T69 = release_idx == 3'h6;
  assign T241 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T70 = T71;
  assign T71 = {T73, T72};
  assign T72 = 2'h0;
  assign T73 = T235;
  assign T74 = T45;
  assign T75 = T76;
  assign T76 = {T78, T77};
  assign T77 = 2'h2;
  assign T78 = 2'h0;
  assign T79 = io_inner_release_valid & T80;
  assign T80 = release_idx == 3'h5;
  assign T242 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T81 = T82;
  assign T82 = {T84, T83};
  assign T83 = 2'h0;
  assign T84 = T235;
  assign T85 = T45;
  assign T86 = T87;
  assign T87 = {T89, T88};
  assign T88 = 2'h2;
  assign T89 = 2'h0;
  assign T90 = io_inner_release_valid & T91;
  assign T91 = release_idx == 3'h4;
  assign T243 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T92 = T93;
  assign T93 = {T95, T94};
  assign T94 = 2'h0;
  assign T95 = T235;
  assign T96 = T45;
  assign T97 = T98;
  assign T98 = {T100, T99};
  assign T99 = 2'h2;
  assign T100 = 2'h0;
  assign T101 = io_inner_release_valid & T102;
  assign T102 = release_idx == 3'h3;
  assign T244 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T103 = T104;
  assign T104 = {T106, T105};
  assign T105 = 2'h0;
  assign T106 = T235;
  assign T107 = T45;
  assign T108 = T109;
  assign T109 = {T111, T110};
  assign T110 = 2'h2;
  assign T111 = 2'h0;
  assign T112 = io_inner_release_valid & T113;
  assign T113 = release_idx == 3'h2;
  assign T245 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T114 = T115;
  assign T115 = {T117, T116};
  assign T116 = 2'h0;
  assign T117 = T235;
  assign T118 = T45;
  assign T119 = T120;
  assign T120 = {T122, T121};
  assign T121 = 2'h2;
  assign T122 = 2'h0;
  assign T123 = io_inner_release_valid & T124;
  assign T124 = release_idx == 3'h1;
  assign T246 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T125 = T126;
  assign T126 = {T128, T127};
  assign T127 = 2'h0;
  assign T128 = T235;
  assign T129 = T45;
  assign T130 = T131;
  assign T131 = {T133, T132};
  assign T132 = 2'h1;
  assign T133 = rel_data_cnt;
  assign T247 = reset ? 2'h0 : T134;
  assign T134 = vwbdq_enq ? T135 : rel_data_cnt;
  assign T135 = rel_data_cnt + 2'h1;
  assign vwbdq_enq = T143 & T136;
  assign T136 = T138 | T137;
  assign T137 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T138 = T140 | T139;
  assign T139 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T140 = T142 | T141;
  assign T141 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T142 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T143 = T144 & voluntary;
  assign voluntary = io_inner_release_bits_payload_r_type == 3'h0;
  assign T144 = io_inner_release_ready & io_inner_release_valid;
  assign T145 = io_inner_release_valid & T146;
  assign T146 = release_idx == 3'h0;
  assign T248 = io_inner_acquire_bits_payload_subblock[4'h9:1'h0];
  assign T147 = T148;
  assign T148 = {T150, T149};
  assign T149 = 2'h0;
  assign T150 = T235;
  assign io_outer_finish_bits_payload_manager_xact_id = outer_arb_io_out_finish_bits_payload_manager_xact_id;
  assign io_outer_finish_bits_header_dst = outer_arb_io_out_finish_bits_header_dst;
  assign io_outer_finish_bits_header_src = outer_arb_io_out_finish_bits_header_src;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_payload_subblock = T249;
  assign T249 = {119'h0, outer_arb_io_out_acquire_bits_payload_subblock};
  assign io_outer_acquire_bits_payload_a_type = outer_arb_io_out_acquire_bits_payload_a_type;
  assign io_outer_acquire_bits_payload_uncached = outer_arb_io_out_acquire_bits_payload_uncached;
  assign io_outer_acquire_bits_payload_data = T151;
  assign T151 = T196 ? T175 : T152;
  assign T152 = T174 ? T153 : io_inner_release_bits_payload_data;
  assign T153 = T173 ? T165 : T154;
  assign T154 = T163 ? vwbdq_1 : vwbdq_0;
  assign T155 = T156 ? io_inner_release_bits_payload_data : vwbdq_0;
  assign T156 = vwbdq_enq & T157;
  assign T157 = T158[1'h0:1'h0];
  assign T158 = 1'h1 << T159;
  assign T159 = rel_data_cnt;
  assign T160 = T161 ? io_inner_release_bits_payload_data : vwbdq_1;
  assign T161 = vwbdq_enq & T162;
  assign T162 = T158[1'h1:1'h1];
  assign T163 = T164[1'h0:1'h0];
  assign T164 = T42;
  assign T165 = T172 ? vwbdq_3 : vwbdq_2;
  assign T166 = T167 ? io_inner_release_bits_payload_data : vwbdq_2;
  assign T167 = vwbdq_enq & T168;
  assign T168 = T158[2'h2:2'h2];
  assign T169 = T170 ? io_inner_release_bits_payload_data : vwbdq_3;
  assign T170 = vwbdq_enq & T171;
  assign T171 = T158[2'h3:2'h3];
  assign T172 = T164[1'h0:1'h0];
  assign T173 = T164[1'h1:1'h1];
  assign T174 = T34 == 2'h1;
  assign T175 = T195 ? T187 : T176;
  assign T176 = T185 ? sdq_1 : sdq_0;
  assign T177 = T178 ? io_inner_acquire_bits_payload_data : sdq_0;
  assign T178 = sdq_enq & T179;
  assign T179 = T180[1'h0:1'h0];
  assign T180 = 1'h1 << T181;
  assign T181 = T235;
  assign T182 = T183 ? io_inner_acquire_bits_payload_data : sdq_1;
  assign T183 = sdq_enq & T184;
  assign T184 = T180[1'h1:1'h1];
  assign T185 = T186[1'h0:1'h0];
  assign T186 = T42;
  assign T187 = T194 ? sdq_3 : sdq_2;
  assign T188 = T189 ? io_inner_acquire_bits_payload_data : sdq_2;
  assign T189 = sdq_enq & T190;
  assign T190 = T180[2'h2:2'h2];
  assign T191 = T192 ? io_inner_acquire_bits_payload_data : sdq_3;
  assign T192 = sdq_enq & T193;
  assign T193 = T180[2'h3:2'h3];
  assign T194 = T186[1'h0:1'h0];
  assign T195 = T186[1'h1:1'h1];
  assign T196 = T34 == 2'h0;
  assign io_outer_acquire_bits_payload_client_xact_id = outer_arb_io_out_acquire_bits_payload_client_xact_id;
  assign io_outer_acquire_bits_payload_addr = outer_arb_io_out_acquire_bits_payload_addr;
  assign io_outer_acquire_bits_header_dst = outer_arb_io_out_acquire_bits_header_dst;
  assign io_outer_acquire_bits_header_src = outer_arb_io_out_acquire_bits_header_src;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T197;
  assign T197 = T211 ? T205 : T198;
  assign T198 = T204 ? T202 : T199;
  assign T199 = T200 ? AcquireTracker_0_io_inner_release_ready : VoluntaryReleaseTracker_io_inner_release_ready;
  assign T200 = T201[1'h0:1'h0];
  assign T201 = release_idx;
  assign T202 = T203 ? AcquireTracker_2_io_inner_release_ready : AcquireTracker_1_io_inner_release_ready;
  assign T203 = T201[1'h0:1'h0];
  assign T204 = T201[1'h1:1'h1];
  assign T205 = T210 ? T208 : T206;
  assign T206 = T207 ? AcquireTracker_4_io_inner_release_ready : AcquireTracker_3_io_inner_release_ready;
  assign T207 = T201[1'h0:1'h0];
  assign T208 = T209 ? AcquireTracker_6_io_inner_release_ready : AcquireTracker_5_io_inner_release_ready;
  assign T209 = T201[1'h0:1'h0];
  assign T210 = T201[1'h1:1'h1];
  assign T211 = T201[2'h2:2'h2];
  assign io_inner_probe_bits_payload_p_type = probe_arb_io_out_bits_payload_p_type;
  assign io_inner_probe_bits_payload_addr = probe_arb_io_out_bits_payload_addr;
  assign io_inner_probe_bits_header_dst = probe_arb_io_out_bits_header_dst;
  assign io_inner_probe_bits_header_src = probe_arb_io_out_bits_header_src;
  assign io_inner_probe_valid = probe_arb_io_out_valid;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_grant_bits_payload_g_type = grant_arb_io_out_bits_payload_g_type;
  assign io_inner_grant_bits_payload_uncached = grant_arb_io_out_bits_payload_uncached;
  assign io_inner_grant_bits_payload_manager_xact_id = grant_arb_io_out_bits_payload_manager_xact_id;
  assign io_inner_grant_bits_payload_client_xact_id = grant_arb_io_out_bits_payload_client_xact_id;
  assign io_inner_grant_bits_payload_data = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = grant_arb_io_out_bits_header_dst;
  assign io_inner_grant_bits_header_src = grant_arb_io_out_bits_header_src;
  assign io_inner_grant_valid = grant_arb_io_out_valid;
  assign io_inner_acquire_ready = T212;
  assign T212 = T214 & T213;
  assign T213 = any_acquire_conflict ^ 1'h1;
  assign T214 = T215 & sdq_rdy;
  assign T215 = T216 | AcquireTracker_6_io_inner_acquire_ready;
  assign T216 = T217 | AcquireTracker_5_io_inner_acquire_ready;
  assign T217 = T218 | AcquireTracker_4_io_inner_acquire_ready;
  assign T218 = T219 | AcquireTracker_3_io_inner_acquire_ready;
  assign T219 = T220 | AcquireTracker_2_io_inner_acquire_ready;
  assign T220 = T221 | AcquireTracker_1_io_inner_acquire_ready;
  assign T221 = VoluntaryReleaseTracker_io_inner_acquire_ready | AcquireTracker_0_io_inner_acquire_ready;
  VoluntaryReleaseTracker VoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_0_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T147 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T248 ),
       .io_inner_grant_ready( grant_arb_io_in_0_ready ),
       .io_inner_grant_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( VoluntaryReleaseTracker_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_0_ready ),
       .io_inner_probe_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_header_src(  )
       //.io_inner_probe_bits_header_dst(  )
       //.io_inner_probe_bits_payload_addr(  )
       //.io_inner_probe_bits_payload_p_type(  )
       .io_inner_release_ready( VoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T145 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T130 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_0_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_0_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T129 ),
       .io_has_acquire_conflict( VoluntaryReleaseTracker_io_has_acquire_conflict ),
       .io_has_release_match( VoluntaryReleaseTracker_io_has_release_match )
  );
  AcquireTracker_0 AcquireTracker_0(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_0_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_1_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T125 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T246 ),
       .io_inner_grant_ready( grant_arb_io_in_1_ready ),
       .io_inner_grant_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_0_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_1_ready ),
       .io_inner_probe_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_0_io_inner_release_ready ),
       .io_inner_release_valid( T123 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T119 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_0_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_0_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_1_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_1_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T118 ),
       .io_has_acquire_conflict( AcquireTracker_0_io_has_acquire_conflict ),
       .io_has_release_match( AcquireTracker_0_io_has_release_match )
  );
  AcquireTracker_1 AcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_2_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T114 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T245 ),
       .io_inner_grant_ready( grant_arb_io_in_2_ready ),
       .io_inner_grant_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_1_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_2_ready ),
       .io_inner_probe_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T112 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T108 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_1_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_1_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_2_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_2_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T107 ),
       .io_has_acquire_conflict( AcquireTracker_1_io_has_acquire_conflict ),
       .io_has_release_match( AcquireTracker_1_io_has_release_match )
  );
  AcquireTracker_2 AcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_3_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T103 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T244 ),
       .io_inner_grant_ready( grant_arb_io_in_3_ready ),
       .io_inner_grant_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_2_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_3_ready ),
       .io_inner_probe_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T101 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T97 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_2_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_2_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_3_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_3_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T96 ),
       .io_has_acquire_conflict( AcquireTracker_2_io_has_acquire_conflict ),
       .io_has_release_match( AcquireTracker_2_io_has_release_match )
  );
  AcquireTracker_3 AcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_4_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T92 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T243 ),
       .io_inner_grant_ready( grant_arb_io_in_4_ready ),
       .io_inner_grant_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_3_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_4_ready ),
       .io_inner_probe_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T90 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T86 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_3_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_3_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_4_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_4_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T85 ),
       .io_has_acquire_conflict( AcquireTracker_3_io_has_acquire_conflict ),
       .io_has_release_match( AcquireTracker_3_io_has_release_match )
  );
  AcquireTracker_4 AcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_5_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T81 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T242 ),
       .io_inner_grant_ready( grant_arb_io_in_5_ready ),
       .io_inner_grant_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_4_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_5_ready ),
       .io_inner_probe_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( T79 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T75 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_4_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_4_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_5_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_5_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T74 ),
       .io_has_acquire_conflict( AcquireTracker_4_io_has_acquire_conflict ),
       .io_has_release_match( AcquireTracker_4_io_has_release_match )
  );
  AcquireTracker_5 AcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_6_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T70 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T241 ),
       .io_inner_grant_ready( grant_arb_io_in_6_ready ),
       .io_inner_grant_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_5_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_6_ready ),
       .io_inner_probe_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( T68 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T64 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_5_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_5_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_6_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_6_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T63 ),
       .io_has_acquire_conflict( AcquireTracker_5_io_has_acquire_conflict ),
       .io_has_release_match( AcquireTracker_5_io_has_release_match )
  );
  AcquireTracker_6 AcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_7_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( T58 ),
       .io_inner_acquire_bits_payload_uncached( io_inner_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( T234 ),
       .io_inner_grant_ready( grant_arb_io_in_7_ready ),
       .io_inner_grant_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( AcquireTracker_6_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( io_inner_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_7_ready ),
       .io_inner_probe_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( T50 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( T46 ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       //.io_outer_acquire_bits_header_src(  )
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( AcquireTracker_6_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( AcquireTracker_6_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( outer_arb_io_in_7_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( outer_arb_io_in_7_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_manager_xact_id(  )
       .io_tile_incoherent( T44 ),
       .io_has_acquire_conflict( AcquireTracker_6_io_has_acquire_conflict )
       //.io_has_release_match(  )
  );
  Arbiter_9 alloc_arb(
       .io_in_7_ready( alloc_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_acquire_ready ),
       //.io_in_7_bits(  )
       .io_in_6_ready( alloc_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_acquire_ready ),
       //.io_in_6_bits(  )
       .io_in_5_ready( alloc_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_acquire_ready ),
       //.io_in_5_bits(  )
       .io_in_4_ready( alloc_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_acquire_ready ),
       //.io_in_4_bits(  )
       .io_in_3_ready( alloc_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_acquire_ready ),
       //.io_in_3_bits(  )
       .io_in_2_ready( alloc_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_acquire_ready ),
       //.io_in_2_bits(  )
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_acquire_ready ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T0 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign alloc_arb.io_in_7_bits = {1{$random}};
    assign alloc_arb.io_in_6_bits = {1{$random}};
    assign alloc_arb.io_in_5_bits = {1{$random}};
    assign alloc_arb.io_in_4_bits = {1{$random}};
    assign alloc_arb.io_in_3_bits = {1{$random}};
    assign alloc_arb.io_in_2_bits = {1{$random}};
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_10 probe_arb(
       .io_in_7_ready( probe_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_in_7_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_in_7_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_in_6_ready( probe_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_in_6_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_in_6_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_in_5_ready( probe_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_in_5_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_in_5_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_in_4_ready( probe_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_in_4_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_in_4_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_in_3_ready( probe_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_in_3_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_in_3_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_in_2_ready( probe_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_in_2_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_in_2_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_in_1_ready( probe_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_in_1_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_in_1_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_in_0_ready( probe_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_p_type(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( probe_arb_io_out_valid ),
       .io_out_bits_header_src( probe_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( probe_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( probe_arb_io_out_bits_payload_addr ),
       .io_out_bits_payload_p_type( probe_arb_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign probe_arb.io_in_0_bits_header_src = {1{$random}};
    assign probe_arb.io_in_0_bits_header_dst = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_addr = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_p_type = {1{$random}};
// synthesis translate_on
`endif
  LockingArbiter_2 grant_arb(.clk(clk), .reset(reset),
       .io_in_7_ready( grant_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_in_7_bits_payload_data( T230 ),
       .io_in_7_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_manager_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_7_bits_payload_uncached( AcquireTracker_6_io_inner_grant_bits_payload_uncached ),
       .io_in_7_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       .io_in_6_ready( grant_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_in_6_bits_payload_data( T229 ),
       .io_in_6_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_manager_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_6_bits_payload_uncached( AcquireTracker_5_io_inner_grant_bits_payload_uncached ),
       .io_in_6_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       .io_in_5_ready( grant_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_in_5_bits_payload_data( T228 ),
       .io_in_5_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_manager_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_5_bits_payload_uncached( AcquireTracker_4_io_inner_grant_bits_payload_uncached ),
       .io_in_5_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       .io_in_4_ready( grant_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_in_4_bits_payload_data( T227 ),
       .io_in_4_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_manager_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_4_bits_payload_uncached( AcquireTracker_3_io_inner_grant_bits_payload_uncached ),
       .io_in_4_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       .io_in_3_ready( grant_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_in_3_bits_payload_data( T226 ),
       .io_in_3_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_manager_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_3_bits_payload_uncached( AcquireTracker_2_io_inner_grant_bits_payload_uncached ),
       .io_in_3_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       .io_in_2_ready( grant_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_in_2_bits_payload_data( T225 ),
       .io_in_2_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_manager_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_2_bits_payload_uncached( AcquireTracker_1_io_inner_grant_bits_payload_uncached ),
       .io_in_2_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       .io_in_1_ready( grant_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_in_1_bits_payload_data( T224 ),
       .io_in_1_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_manager_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_1_bits_payload_uncached( AcquireTracker_0_io_inner_grant_bits_payload_uncached ),
       .io_in_1_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       .io_in_0_ready( grant_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_in_0_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_in_0_bits_payload_data( T223 ),
       .io_in_0_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_uncached( VoluntaryReleaseTracker_io_inner_grant_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( grant_arb_io_out_valid ),
       .io_out_bits_header_src( grant_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( grant_arb_io_out_bits_header_dst ),
       //.io_out_bits_payload_data(  )
       .io_out_bits_payload_client_xact_id( grant_arb_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( grant_arb_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( grant_arb_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( grant_arb_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  UncachedTileLinkIOArbiterThatPassesId outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       //.io_in_7_acquire_bits_header_src(  )
       //.io_in_7_acquire_bits_header_dst(  )
       .io_in_7_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_in_7_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_7_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_in_7_acquire_bits_payload_uncached( AcquireTracker_6_io_outer_acquire_bits_payload_uncached ),
       .io_in_7_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_in_7_acquire_bits_payload_subblock( AcquireTracker_6_io_outer_acquire_bits_payload_subblock ),
       .io_in_7_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_in_7_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_in_7_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_in_7_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_in_7_grant_bits_payload_manager_xact_id( outer_arb_io_in_7_grant_bits_payload_manager_xact_id ),
       .io_in_7_grant_bits_payload_uncached( outer_arb_io_in_7_grant_bits_payload_uncached ),
       .io_in_7_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_in_7_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_in_7_finish_valid(  )
       //.io_in_7_finish_bits_header_src(  )
       //.io_in_7_finish_bits_header_dst(  )
       //.io_in_7_finish_bits_payload_manager_xact_id(  )
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       //.io_in_6_acquire_bits_header_src(  )
       //.io_in_6_acquire_bits_header_dst(  )
       .io_in_6_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_in_6_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_6_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_in_6_acquire_bits_payload_uncached( AcquireTracker_5_io_outer_acquire_bits_payload_uncached ),
       .io_in_6_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_in_6_acquire_bits_payload_subblock( AcquireTracker_5_io_outer_acquire_bits_payload_subblock ),
       .io_in_6_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_in_6_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_in_6_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_in_6_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_in_6_grant_bits_payload_manager_xact_id( outer_arb_io_in_6_grant_bits_payload_manager_xact_id ),
       .io_in_6_grant_bits_payload_uncached( outer_arb_io_in_6_grant_bits_payload_uncached ),
       .io_in_6_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_in_6_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_in_6_finish_valid(  )
       //.io_in_6_finish_bits_header_src(  )
       //.io_in_6_finish_bits_header_dst(  )
       //.io_in_6_finish_bits_payload_manager_xact_id(  )
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       //.io_in_5_acquire_bits_header_src(  )
       //.io_in_5_acquire_bits_header_dst(  )
       .io_in_5_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_in_5_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_5_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_in_5_acquire_bits_payload_uncached( AcquireTracker_4_io_outer_acquire_bits_payload_uncached ),
       .io_in_5_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_in_5_acquire_bits_payload_subblock( AcquireTracker_4_io_outer_acquire_bits_payload_subblock ),
       .io_in_5_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_in_5_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_in_5_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_in_5_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_in_5_grant_bits_payload_manager_xact_id( outer_arb_io_in_5_grant_bits_payload_manager_xact_id ),
       .io_in_5_grant_bits_payload_uncached( outer_arb_io_in_5_grant_bits_payload_uncached ),
       .io_in_5_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_in_5_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_in_5_finish_valid(  )
       //.io_in_5_finish_bits_header_src(  )
       //.io_in_5_finish_bits_header_dst(  )
       //.io_in_5_finish_bits_payload_manager_xact_id(  )
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       //.io_in_4_acquire_bits_header_src(  )
       //.io_in_4_acquire_bits_header_dst(  )
       .io_in_4_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_in_4_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_4_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_in_4_acquire_bits_payload_uncached( AcquireTracker_3_io_outer_acquire_bits_payload_uncached ),
       .io_in_4_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_in_4_acquire_bits_payload_subblock( AcquireTracker_3_io_outer_acquire_bits_payload_subblock ),
       .io_in_4_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_in_4_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_in_4_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_in_4_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_in_4_grant_bits_payload_manager_xact_id( outer_arb_io_in_4_grant_bits_payload_manager_xact_id ),
       .io_in_4_grant_bits_payload_uncached( outer_arb_io_in_4_grant_bits_payload_uncached ),
       .io_in_4_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_in_4_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_in_4_finish_valid(  )
       //.io_in_4_finish_bits_header_src(  )
       //.io_in_4_finish_bits_header_dst(  )
       //.io_in_4_finish_bits_payload_manager_xact_id(  )
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       //.io_in_3_acquire_bits_header_src(  )
       //.io_in_3_acquire_bits_header_dst(  )
       .io_in_3_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_in_3_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_3_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_in_3_acquire_bits_payload_uncached( AcquireTracker_2_io_outer_acquire_bits_payload_uncached ),
       .io_in_3_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_in_3_acquire_bits_payload_subblock( AcquireTracker_2_io_outer_acquire_bits_payload_subblock ),
       .io_in_3_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_in_3_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_in_3_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_in_3_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_in_3_grant_bits_payload_manager_xact_id( outer_arb_io_in_3_grant_bits_payload_manager_xact_id ),
       .io_in_3_grant_bits_payload_uncached( outer_arb_io_in_3_grant_bits_payload_uncached ),
       .io_in_3_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_in_3_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_in_3_finish_valid(  )
       //.io_in_3_finish_bits_header_src(  )
       //.io_in_3_finish_bits_header_dst(  )
       //.io_in_3_finish_bits_payload_manager_xact_id(  )
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       //.io_in_2_acquire_bits_header_src(  )
       //.io_in_2_acquire_bits_header_dst(  )
       .io_in_2_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_uncached( AcquireTracker_1_io_outer_acquire_bits_payload_uncached ),
       .io_in_2_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_subblock( AcquireTracker_1_io_outer_acquire_bits_payload_subblock ),
       .io_in_2_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_manager_xact_id( outer_arb_io_in_2_grant_bits_payload_manager_xact_id ),
       .io_in_2_grant_bits_payload_uncached( outer_arb_io_in_2_grant_bits_payload_uncached ),
       .io_in_2_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_in_2_finish_valid(  )
       //.io_in_2_finish_bits_header_src(  )
       //.io_in_2_finish_bits_header_dst(  )
       //.io_in_2_finish_bits_payload_manager_xact_id(  )
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       //.io_in_1_acquire_bits_header_src(  )
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_uncached( AcquireTracker_0_io_outer_acquire_bits_payload_uncached ),
       .io_in_1_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_subblock( AcquireTracker_0_io_outer_acquire_bits_payload_subblock ),
       .io_in_1_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_manager_xact_id( outer_arb_io_in_1_grant_bits_payload_manager_xact_id ),
       .io_in_1_grant_bits_payload_uncached( outer_arb_io_in_1_grant_bits_payload_uncached ),
       .io_in_1_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_in_1_finish_valid(  )
       //.io_in_1_finish_bits_header_src(  )
       //.io_in_1_finish_bits_header_dst(  )
       //.io_in_1_finish_bits_payload_manager_xact_id(  )
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       //.io_in_0_acquire_bits_header_src(  )
       //.io_in_0_acquire_bits_header_dst(  )
       .io_in_0_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_uncached( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_uncached ),
       .io_in_0_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_subblock( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subblock ),
       .io_in_0_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_manager_xact_id( outer_arb_io_in_0_grant_bits_payload_manager_xact_id ),
       .io_in_0_grant_bits_payload_uncached( outer_arb_io_in_0_grant_bits_payload_uncached ),
       .io_in_0_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_in_0_finish_valid(  )
       //.io_in_0_finish_bits_header_src(  )
       //.io_in_0_finish_bits_header_dst(  )
       //.io_in_0_finish_bits_payload_manager_xact_id(  )
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( outer_arb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( outer_arb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( outer_arb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( outer_arb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( outer_arb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_uncached( outer_arb_io_out_acquire_bits_payload_uncached ),
       .io_out_acquire_bits_payload_a_type( outer_arb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_subblock( outer_arb_io_out_acquire_bits_payload_subblock ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_header_src( io_outer_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_outer_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( T222 ),
       .io_out_grant_bits_payload_client_xact_id( io_outer_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_manager_xact_id( io_outer_grant_bits_payload_manager_xact_id ),
       .io_out_grant_bits_payload_uncached( io_outer_grant_bits_payload_uncached ),
       .io_out_grant_bits_payload_g_type( io_outer_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_outer_finish_ready ),
       .io_out_finish_valid( outer_arb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( outer_arb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( outer_arb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_manager_xact_id( outer_arb_io_out_finish_bits_payload_manager_xact_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign outer_arb.io_in_7_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_7_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_valid = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_6_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_6_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_valid = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_5_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_5_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_valid = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_4_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_valid = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_valid = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_valid = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_valid = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_payload_manager_xact_id = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_valid = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_payload_manager_xact_id = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      sdq_val <= 4'h0;
    end else if(T43) begin
      sdq_val <= T11;
    end
    if(reset) begin
      rel_data_cnt <= 2'h0;
    end else if(vwbdq_enq) begin
      rel_data_cnt <= T135;
    end
    if(T156) begin
      vwbdq_0 <= io_inner_release_bits_payload_data;
    end
    if(T161) begin
      vwbdq_1 <= io_inner_release_bits_payload_data;
    end
    if(T167) begin
      vwbdq_2 <= io_inner_release_bits_payload_data;
    end
    if(T170) begin
      vwbdq_3 <= io_inner_release_bits_payload_data;
    end
    if(T178) begin
      sdq_0 <= io_inner_acquire_bits_payload_data;
    end
    if(T183) begin
      sdq_1 <= io_inner_acquire_bits_payload_data;
    end
    if(T189) begin
      sdq_2 <= io_inner_acquire_bits_payload_data;
    end
    if(T192) begin
      sdq_3 <= io_inner_acquire_bits_payload_data;
    end
  end
endmodule

module TagCacheMetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_id,
    input [16:0] io_read_bits_tag,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [16:0] io_write_bits_tag,
    input [5:0] io_write_bits_idx,
    input [7:0] io_write_bits_way_en,
    output io_resp_valid,
    output io_resp_bits_id,
    output[16:0] io_resp_bits_tag,
    output io_resp_bits_hit,
    output[7:0] io_resp_bits_way_en
);

  wire[7:0] T0;
  reg [7:0] s2_replace_way;
  wire[7:0] T1;
  wire[7:0] s1_replace_way;
  wire[2:0] T2;
  reg [15:0] R3;
  wire[15:0] T99;
  wire[15:0] T4;
  wire[15:0] T5;
  wire[14:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  s1_clk_en;
  wire T15;
  reg [7:0] s2_match_way;
  wire[7:0] T16;
  wire[7:0] s1_match_way;
  wire[7:0] T17;
  wire[3:0] T18;
  wire[1:0] T19;
  wire T20;
  reg [16:0] s1_tag;
  wire[16:0] T21;
  wire[16:0] T22;
  wire[135:0] ctags;
  wire[135:0] T23;
  wire[135:0] T24;
  wire[135:0] T25;
  wire[67:0] T26;
  wire[33:0] T27;
  wire[16:0] T28;
  wire[16:0] T100;
  wire T29;
  wire[7:0] wmask;
  wire rst;
  reg [6:0] rst_cnt;
  wire[6:0] T101;
  wire[6:0] T30;
  wire[6:0] T31;
  wire[16:0] T32;
  wire[16:0] T102;
  wire T33;
  wire[33:0] T34;
  wire[16:0] T35;
  wire[16:0] T103;
  wire T36;
  wire[16:0] T37;
  wire[16:0] T104;
  wire T38;
  wire[67:0] T39;
  wire[33:0] T40;
  wire[16:0] T41;
  wire[16:0] T105;
  wire T42;
  wire[16:0] T43;
  wire[16:0] T106;
  wire T44;
  wire[33:0] T45;
  wire[16:0] T46;
  wire[16:0] T107;
  wire T47;
  wire[16:0] T48;
  wire[16:0] T108;
  wire T49;
  wire[135:0] T50;
  wire[67:0] T51;
  wire[33:0] T52;
  wire[16:0] wdata;
  wire T53;
  wire[5:0] T109;
  wire[6:0] waddr;
  wire[6:0] T110;
  reg [5:0] R54;
  wire[5:0] T55;
  wire T56;
  wire[16:0] T57;
  wire[1:0] T58;
  wire T59;
  wire[16:0] T60;
  wire T61;
  wire[16:0] T62;
  wire[3:0] T63;
  wire[1:0] T64;
  wire T65;
  wire[16:0] T66;
  wire T67;
  wire[16:0] T68;
  wire[1:0] T69;
  wire T70;
  wire[16:0] T71;
  wire T72;
  wire[16:0] T73;
  reg  s2_hit;
  wire T74;
  wire s1_hit;
  reg [16:0] s2_replace_meta;
  wire[16:0] T75;
  wire[16:0] s1_replace_meta;
  wire[16:0] T76;
  wire[16:0] T77;
  wire T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[16:0] T81;
  wire T82;
  wire T83;
  wire[16:0] T84;
  wire[16:0] T85;
  wire T86;
  wire[16:0] T87;
  wire T88;
  wire T89;
  wire T90;
  reg  R91;
  wire T92;
  reg  s1_id;
  wire T93;
  reg  R94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s2_replace_way = {1{$random}};
    R3 = {1{$random}};
    s1_clk_en = {1{$random}};
    s2_match_way = {1{$random}};
    s1_tag = {1{$random}};
    rst_cnt = {1{$random}};
    R54 = {1{$random}};
    s2_hit = {1{$random}};
    s2_replace_meta = {1{$random}};
    R91 = {1{$random}};
    s1_id = {1{$random}};
    R94 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_way_en = T0;
  assign T0 = s2_hit ? s2_match_way : s2_replace_way;
  assign T1 = s1_clk_en ? s1_replace_way : s2_replace_way;
  assign s1_replace_way = 1'h1 << T2;
  assign T2 = R3[2'h2:1'h0];
  assign T99 = reset ? 16'h1 : T4;
  assign T4 = T14 ? T5 : R3;
  assign T5 = {T7, T6};
  assign T6 = R3[4'hf:1'h1];
  assign T7 = T9 ^ T8;
  assign T8 = R3[3'h5:3'h5];
  assign T9 = T11 ^ T10;
  assign T10 = R3[2'h3:2'h3];
  assign T11 = T13 ^ T12;
  assign T12 = R3[2'h2:2'h2];
  assign T13 = R3[1'h0:1'h0];
  assign T14 = 1'h0;
  assign T15 = io_read_ready & io_read_valid;
  assign T16 = s1_clk_en ? s1_match_way : s2_match_way;
  assign s1_match_way = T17;
  assign T17 = {T63, T18};
  assign T18 = {T58, T19};
  assign T19 = {T56, T20};
  assign T20 = T22 == s1_tag;
  assign T21 = io_read_valid ? io_read_bits_tag : s1_tag;
  assign T22 = ctags[5'h10:1'h0];
  TagCacheMetadataArray_metaArray metaArray (
    .CLK(clk),
    .W0A(T109),
    .W0E(T53),
    .W0I(T50),
    .W0M(T24),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(ctags)
  );
  assign T24 = T25;
  assign T25 = {T39, T26};
  assign T26 = {T34, T27};
  assign T27 = {T32, T28};
  assign T28 = 17'h0 - T100;
  assign T100 = {16'h0, T29};
  assign T29 = wmask[1'h0:1'h0];
  assign wmask = rst ? 8'hff : io_write_bits_way_en;
  assign rst = rst_cnt < 7'h40;
  assign T101 = reset ? 7'h0 : T30;
  assign T30 = rst ? T31 : rst_cnt;
  assign T31 = rst_cnt + 7'h1;
  assign T32 = 17'h0 - T102;
  assign T102 = {16'h0, T33};
  assign T33 = wmask[1'h1:1'h1];
  assign T34 = {T37, T35};
  assign T35 = 17'h0 - T103;
  assign T103 = {16'h0, T36};
  assign T36 = wmask[2'h2:2'h2];
  assign T37 = 17'h0 - T104;
  assign T104 = {16'h0, T38};
  assign T38 = wmask[2'h3:2'h3];
  assign T39 = {T45, T40};
  assign T40 = {T43, T41};
  assign T41 = 17'h0 - T105;
  assign T105 = {16'h0, T42};
  assign T42 = wmask[3'h4:3'h4];
  assign T43 = 17'h0 - T106;
  assign T106 = {16'h0, T44};
  assign T44 = wmask[3'h5:3'h5];
  assign T45 = {T48, T46};
  assign T46 = 17'h0 - T107;
  assign T107 = {16'h0, T47};
  assign T47 = wmask[3'h6:3'h6];
  assign T48 = 17'h0 - T108;
  assign T108 = {16'h0, T49};
  assign T49 = wmask[3'h7:3'h7];
  assign T50 = {T51, T51};
  assign T51 = {T52, T52};
  assign T52 = {wdata, wdata};
  assign wdata = rst ? 17'h0 : io_write_bits_tag;
  assign T53 = rst | io_write_valid;
  assign T109 = waddr[3'h5:1'h0];
  assign waddr = rst ? rst_cnt : T110;
  assign T110 = {1'h0, io_write_bits_idx};
  assign T55 = io_read_valid ? io_read_bits_idx : R54;
  assign T56 = T57 == s1_tag;
  assign T57 = ctags[6'h21:5'h11];
  assign T58 = {T61, T59};
  assign T59 = T60 == s1_tag;
  assign T60 = ctags[6'h32:6'h22];
  assign T61 = T62 == s1_tag;
  assign T62 = ctags[7'h43:6'h33];
  assign T63 = {T69, T64};
  assign T64 = {T67, T65};
  assign T65 = T66 == s1_tag;
  assign T66 = ctags[7'h54:7'h44];
  assign T67 = T68 == s1_tag;
  assign T68 = ctags[7'h65:7'h55];
  assign T69 = {T72, T70};
  assign T70 = T71 == s1_tag;
  assign T71 = ctags[7'h76:7'h66];
  assign T72 = T73 == s1_tag;
  assign T73 = ctags[8'h87:7'h77];
  assign T74 = s1_clk_en ? s1_hit : s2_hit;
  assign s1_hit = s1_match_way != 8'h0;
  assign io_resp_bits_hit = s2_hit;
  assign io_resp_bits_tag = s2_replace_meta;
  assign T75 = s1_clk_en ? s1_replace_meta : s2_replace_meta;
  assign s1_replace_meta = T90 ? T84 : T76;
  assign T76 = T83 ? T81 : T77;
  assign T77 = T78 ? T57 : T22;
  assign T78 = T79[1'h0:1'h0];
  assign T79 = T80;
  assign T80 = R3[2'h2:1'h0];
  assign T81 = T82 ? T62 : T60;
  assign T82 = T79[1'h0:1'h0];
  assign T83 = T79[1'h1:1'h1];
  assign T84 = T89 ? T87 : T85;
  assign T85 = T86 ? T68 : T66;
  assign T86 = T79[1'h0:1'h0];
  assign T87 = T88 ? T73 : T71;
  assign T88 = T79[1'h0:1'h0];
  assign T89 = T79[1'h1:1'h1];
  assign T90 = T79[2'h2:2'h2];
  assign io_resp_bits_id = R91;
  assign T92 = s1_clk_en ? s1_id : R91;
  assign T93 = io_read_valid ? io_read_bits_id : s1_id;
  assign io_resp_valid = R94;
  assign io_write_ready = T95;
  assign T95 = rst ^ 1'h1;
  assign io_read_ready = T96;
  assign T96 = T98 & T97;
  assign T97 = io_write_valid ^ 1'h1;
  assign T98 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(s1_clk_en) begin
      s2_replace_way <= s1_replace_way;
    end
    if(reset) begin
      R3 <= 16'h1;
    end else if(T14) begin
      R3 <= T5;
    end
    s1_clk_en <= T15;
    if(s1_clk_en) begin
      s2_match_way <= s1_match_way;
    end
    if(io_read_valid) begin
      s1_tag <= io_read_bits_tag;
    end
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(rst) begin
      rst_cnt <= T31;
    end
    if(io_read_valid) begin
      R54 <= io_read_bits_idx;
    end
    if(s1_clk_en) begin
      s2_hit <= s1_hit;
    end
    if(s1_clk_en) begin
      s2_replace_meta <= s1_replace_meta;
    end
    if(s1_clk_en) begin
      R91 <= s1_id;
    end
    if(io_read_valid) begin
      s1_id <= io_read_bits_id;
    end
    R94 <= s1_clk_en;
  end
endmodule

module TagCacheDataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_id,
    input [7:0] io_read_bits_addr,
    input [7:0] io_read_bits_way_en,
    output io_write_ready,
    input  io_write_valid,
    input [127:0] io_write_bits_data,
    input [7:0] io_write_bits_addr,
    input [7:0] io_write_bits_way_en,
    input [3:0] io_write_bits_wmask,
    output io_resp_valid,
    output io_resp_bits_id,
    output[127:0] io_resp_bits_data
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[127:0] resp_7;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T15;
  wire T16;
  wire[127:0] T3;
  wire[127:0] wmask;
  wire[127:0] T4;
  wire[63:0] T5;
  wire[31:0] T6;
  wire[31:0] T119;
  wire T7;
  wire[31:0] T8;
  wire[31:0] T120;
  wire T9;
  wire[63:0] T10;
  wire[31:0] T11;
  wire[31:0] T121;
  wire T12;
  wire[31:0] T13;
  wire[31:0] T122;
  wire T14;
  reg [7:0] R17;
  wire[7:0] T18;
  wire T23;
  reg [7:0] R24;
  wire[127:0] T25;
  wire[127:0] T26;
  wire[127:0] resp_6;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T29;
  wire T30;
  wire[127:0] T28;
  reg [7:0] R31;
  wire[7:0] T32;
  wire T37;
  wire[127:0] T38;
  wire[127:0] T39;
  wire[127:0] resp_5;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T42;
  wire T43;
  wire[127:0] T41;
  reg [7:0] R44;
  wire[7:0] T45;
  wire T50;
  wire[127:0] T51;
  wire[127:0] T52;
  wire[127:0] resp_4;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T55;
  wire T56;
  wire[127:0] T54;
  reg [7:0] R57;
  wire[7:0] T58;
  wire T63;
  wire[127:0] T64;
  wire[127:0] T65;
  wire[127:0] resp_3;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T68;
  wire T69;
  wire[127:0] T67;
  reg [7:0] R70;
  wire[7:0] T71;
  wire T76;
  wire[127:0] T77;
  wire[127:0] T78;
  wire[127:0] resp_2;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T81;
  wire T82;
  wire[127:0] T80;
  reg [7:0] R83;
  wire[7:0] T84;
  wire T89;
  wire[127:0] T90;
  wire[127:0] T91;
  wire[127:0] resp_1;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T94;
  wire T95;
  wire[127:0] T93;
  reg [7:0] R96;
  wire[7:0] T97;
  wire T102;
  wire[127:0] T103;
  wire[127:0] resp_0;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T106;
  wire T107;
  wire[127:0] T105;
  reg [7:0] R108;
  wire[7:0] T109;
  wire T114;
  reg  R115;
  reg  R116;
  wire T117;
  wire T118;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
    R24 = {1{$random}};
    R31 = {1{$random}};
    R44 = {1{$random}};
    R57 = {1{$random}};
    R70 = {1{$random}};
    R83 = {1{$random}};
    R96 = {1{$random}};
    R108 = {1{$random}};
    R115 = {1{$random}};
    R116 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_data = T0;
  assign T0 = T25 | T1;
  assign T1 = T23 ? resp_7 : 128'h0;
  assign T19 = T22 & T20;
  assign T20 = T21 & io_read_valid;
  assign T21 = io_read_bits_way_en[3'h7:3'h7];
  assign T22 = T15 ^ 1'h1;
  assign T15 = T16 & io_write_valid;
  assign T16 = io_write_bits_way_en[3'h7:3'h7];
  TagCacheDataArray_T2 T2 (
    .CLK(clk),
    .RW0A(T15 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T19 || T15),
    .RW0W(T15),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_7)
  );
  assign wmask = T4;
  assign T4 = {T10, T5};
  assign T5 = {T8, T6};
  assign T6 = 32'h0 - T119;
  assign T119 = {31'h0, T7};
  assign T7 = io_write_bits_wmask[1'h0:1'h0];
  assign T8 = 32'h0 - T120;
  assign T120 = {31'h0, T9};
  assign T9 = io_write_bits_wmask[1'h1:1'h1];
  assign T10 = {T13, T11};
  assign T11 = 32'h0 - T121;
  assign T121 = {31'h0, T12};
  assign T12 = io_write_bits_wmask[2'h2:2'h2];
  assign T13 = 32'h0 - T122;
  assign T122 = {31'h0, T14};
  assign T14 = io_write_bits_wmask[2'h3:2'h3];
  assign T18 = T19 ? io_read_bits_addr : R17;
  assign T23 = R24[3'h7:3'h7];
  assign T25 = T38 | T26;
  assign T26 = T37 ? resp_6 : 128'h0;
  assign T33 = T36 & T34;
  assign T34 = T35 & io_read_valid;
  assign T35 = io_read_bits_way_en[3'h6:3'h6];
  assign T36 = T29 ^ 1'h1;
  assign T29 = T30 & io_write_valid;
  assign T30 = io_write_bits_way_en[3'h6:3'h6];
  TagCacheDataArray_T2 T27 (
    .CLK(clk),
    .RW0A(T29 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T33 || T29),
    .RW0W(T29),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_6)
  );
  assign T32 = T33 ? io_read_bits_addr : R31;
  assign T37 = R24[3'h6:3'h6];
  assign T38 = T51 | T39;
  assign T39 = T50 ? resp_5 : 128'h0;
  assign T46 = T49 & T47;
  assign T47 = T48 & io_read_valid;
  assign T48 = io_read_bits_way_en[3'h5:3'h5];
  assign T49 = T42 ^ 1'h1;
  assign T42 = T43 & io_write_valid;
  assign T43 = io_write_bits_way_en[3'h5:3'h5];
  TagCacheDataArray_T2 T40 (
    .CLK(clk),
    .RW0A(T42 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T46 || T42),
    .RW0W(T42),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_5)
  );
  assign T45 = T46 ? io_read_bits_addr : R44;
  assign T50 = R24[3'h5:3'h5];
  assign T51 = T64 | T52;
  assign T52 = T63 ? resp_4 : 128'h0;
  assign T59 = T62 & T60;
  assign T60 = T61 & io_read_valid;
  assign T61 = io_read_bits_way_en[3'h4:3'h4];
  assign T62 = T55 ^ 1'h1;
  assign T55 = T56 & io_write_valid;
  assign T56 = io_write_bits_way_en[3'h4:3'h4];
  TagCacheDataArray_T2 T53 (
    .CLK(clk),
    .RW0A(T55 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T59 || T55),
    .RW0W(T55),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_4)
  );
  assign T58 = T59 ? io_read_bits_addr : R57;
  assign T63 = R24[3'h4:3'h4];
  assign T64 = T77 | T65;
  assign T65 = T76 ? resp_3 : 128'h0;
  assign T72 = T75 & T73;
  assign T73 = T74 & io_read_valid;
  assign T74 = io_read_bits_way_en[2'h3:2'h3];
  assign T75 = T68 ^ 1'h1;
  assign T68 = T69 & io_write_valid;
  assign T69 = io_write_bits_way_en[2'h3:2'h3];
  TagCacheDataArray_T2 T66 (
    .CLK(clk),
    .RW0A(T68 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T72 || T68),
    .RW0W(T68),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_3)
  );
  assign T71 = T72 ? io_read_bits_addr : R70;
  assign T76 = R24[2'h3:2'h3];
  assign T77 = T90 | T78;
  assign T78 = T89 ? resp_2 : 128'h0;
  assign T85 = T88 & T86;
  assign T86 = T87 & io_read_valid;
  assign T87 = io_read_bits_way_en[2'h2:2'h2];
  assign T88 = T81 ^ 1'h1;
  assign T81 = T82 & io_write_valid;
  assign T82 = io_write_bits_way_en[2'h2:2'h2];
  TagCacheDataArray_T2 T79 (
    .CLK(clk),
    .RW0A(T81 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T85 || T81),
    .RW0W(T81),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_2)
  );
  assign T84 = T85 ? io_read_bits_addr : R83;
  assign T89 = R24[2'h2:2'h2];
  assign T90 = T103 | T91;
  assign T91 = T102 ? resp_1 : 128'h0;
  assign T98 = T101 & T99;
  assign T99 = T100 & io_read_valid;
  assign T100 = io_read_bits_way_en[1'h1:1'h1];
  assign T101 = T94 ^ 1'h1;
  assign T94 = T95 & io_write_valid;
  assign T95 = io_write_bits_way_en[1'h1:1'h1];
  TagCacheDataArray_T2 T92 (
    .CLK(clk),
    .RW0A(T94 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T98 || T94),
    .RW0W(T94),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_1)
  );
  assign T97 = T98 ? io_read_bits_addr : R96;
  assign T102 = R24[1'h1:1'h1];
  assign T103 = T114 ? resp_0 : 128'h0;
  assign T110 = T113 & T111;
  assign T111 = T112 & io_read_valid;
  assign T112 = io_read_bits_way_en[1'h0:1'h0];
  assign T113 = T106 ^ 1'h1;
  assign T106 = T107 & io_write_valid;
  assign T107 = io_write_bits_way_en[1'h0:1'h0];
  TagCacheDataArray_T2 T104 (
    .CLK(clk),
    .RW0A(T106 ? io_write_bits_addr : io_read_bits_addr),
    .RW0E(T110 || T106),
    .RW0W(T106),
    .RW0I(io_write_bits_data),
    .RW0M(wmask),
    .RW0O(resp_0)
  );
  assign T109 = T110 ? io_read_bits_addr : R108;
  assign T114 = R24[1'h0:1'h0];
  assign io_resp_bits_id = R115;
  assign io_resp_valid = R116;
  assign T117 = io_read_ready & io_read_valid;
  assign io_write_ready = 1'h1;
  assign io_read_ready = T118;
  assign T118 = io_write_valid ^ 1'h1;

  always @(posedge clk) begin
    if(T19) begin
      R17 <= io_read_bits_addr;
    end
    R24 <= io_read_bits_way_en;
    if(T33) begin
      R31 <= io_read_bits_addr;
    end
    if(T46) begin
      R44 <= io_read_bits_addr;
    end
    if(T59) begin
      R57 <= io_read_bits_addr;
    end
    if(T72) begin
      R70 <= io_read_bits_addr;
    end
    if(T85) begin
      R83 <= io_read_bits_addr;
    end
    if(T98) begin
      R96 <= io_read_bits_addr;
    end
    if(T110) begin
      R108 <= io_read_bits_addr;
    end
    R115 <= io_read_bits_id;
    R116 <= T117;
  end
endmodule

module TagCacheTracker(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [4:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [135:0] io_uncached_acquire_bits_payload_data,
    input  io_uncached_acquire_bits_payload_uncached,
    input [1:0] io_uncached_acquire_bits_payload_a_type,
    input [128:0] io_uncached_acquire_bits_payload_subblock,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[135:0] io_uncached_grant_bits_payload_data,
    output[4:0] io_uncached_grant_bits_payload_client_xact_id,
    output io_uncached_grant_bits_payload_manager_xact_id,
    output io_uncached_grant_bits_payload_uncached,
    output[1:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    //input  io_uncached_finish_valid
    //input [1:0] io_uncached_finish_bits_header_src
    //input [1:0] io_uncached_finish_bits_header_dst
    //input  io_uncached_finish_bits_payload_manager_xact_id
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output io_meta_read_bits_id,
    output[16:0] io_meta_read_bits_tag,
    output[5:0] io_meta_read_bits_idx,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[16:0] io_meta_write_bits_tag,
    output[5:0] io_meta_write_bits_idx,
    output[7:0] io_meta_write_bits_way_en,
    input  io_meta_resp_valid,
    input  io_meta_resp_bits_id,
    input [16:0] io_meta_resp_bits_tag,
    input  io_meta_resp_bits_hit,
    input [7:0] io_meta_resp_bits_way_en,
    input  io_data_read_ready,
    output io_data_read_valid,
    output io_data_read_bits_id,
    output[7:0] io_data_read_bits_addr,
    output[7:0] io_data_read_bits_way_en,
    input  io_data_write_ready,
    output io_data_write_valid,
    output[127:0] io_data_write_bits_data,
    output[7:0] io_data_write_bits_addr,
    output[7:0] io_data_write_bits_way_en,
    output[3:0] io_data_write_bits_wmask,
    input  io_data_resp_valid,
    input  io_data_resp_bits_id,
    input [127:0] io_data_resp_bits_data,
    output io_acq_conflict,
    output io_acq_match
);

  wire T0;
  reg  collect_acq_data;
  wire T431;
  wire T1;
  wire T2;
  wire T3;
  wire acq_data_done;
  wire T4;
  reg [1:0] acq_data_cnt;
  wire[1:0] T432;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T11;
  wire T12;
  wire T13;
  reg [3:0] state;
  wire[3:0] T433;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire T29;
  wire T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire T33;
  wire[3:0] T34;
  reg  acq_wr;
  wire T434;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire wb_read_done;
  wire T48;
  reg [1:0] wb_read_cnt;
  wire[1:0] T435;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire wb_data_done;
  wire T56;
  reg [1:0] wb_data_cnt;
  wire[1:0] T436;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  reg  mem_tag_cmd_sent;
  wire T437;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  reg  acq_data_process;
  wire T438;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  reg  mem_acq_data_sent;
  wire T439;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire mem_acq_data_write_done;
  wire T79;
  reg [1:0] mem_acq_data_write_cnt;
  wire[1:0] T440;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg  mem_acq_cmd_sent;
  wire T441;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  reg  mem_tag_data_sent;
  wire T442;
  wire T95;
  wire T96;
  wire T97;
  wire mem_tag_data_write_done;
  wire T98;
  reg [1:0] mem_tag_data_write_cnt;
  wire[1:0] T443;
  wire[1:0] T99;
  wire[1:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire refill_data_done;
  wire T112;
  reg [1:0] refill_data_cnt;
  wire[1:0] T444;
  wire[1:0] T113;
  wire[1:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire[3:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  reg  gnt_enable;
  wire T445;
  wire T127;
  wire T128;
  wire T129;
  wire gnt_data_done;
  wire T130;
  reg [1:0] gnt_data_cnt;
  wire[1:0] T446;
  wire[1:0] T131;
  wire[1:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  reg  mem_acq_gnt_ready;
  wire T447;
  wire T137;
  wire T138;
  wire T139;
  wire mem_acq_data_read_done;
  wire T140;
  reg [1:0] mem_acq_data_read_cnt;
  wire[1:0] T448;
  wire[1:0] T141;
  wire[1:0] T142;
  wire T143;
  wire mem_resp_is_acq;
  wire T144;
  wire T145;
  wire T146;
  wire acq_has_data;
  wire T8;
  wire T9;
  wire T10;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  reg [25:0] acq_addr;
  wire[25:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[5:0] T157;
  wire[5:0] T158;
  wire[3:0] T159;
  wire[3:0] T160;
  wire[1:0] T161;
  wire T162;
  reg  mem_tag_refill_ready;
  wire T449;
  wire T163;
  wire T164;
  wire T165;
  wire mem_tag_data_read_done;
  wire T166;
  reg [1:0] mem_tag_data_read_cnt;
  wire[1:0] T450;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire mem_resp_is_tag;
  wire T170;
  wire T171;
  wire T172;
  reg [7:0] acq_way_en;
  wire[7:0] T451;
  wire[7:0] T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire[7:0] T177;
  wire[7:0] T178;
  wire[5:0] T179;
  wire[127:0] T452;
  wire[286:0] T180;
  wire[286:0] T181;
  wire[7:0] T182;
  wire[1:0] T183;
  wire[31:0] T184;
  wire[31:0] T185;
  wire[15:0] T186;
  wire[7:0] T187;
  wire[3:0] T188;
  wire[543:0] T189;
  wire[543:0] T190;
  wire[271:0] T191;
  reg [135:0] acq_data_0;
  wire[135:0] T192;
  wire T193;
  wire T194;
  wire[3:0] T195;
  wire[1:0] T196;
  wire T197;
  reg [135:0] acq_data_1;
  wire[135:0] T198;
  wire T199;
  wire T200;
  wire[271:0] T201;
  reg [135:0] acq_data_2;
  wire[135:0] T202;
  wire T203;
  wire T204;
  reg [135:0] acq_data_3;
  wire[135:0] T205;
  wire T206;
  wire T207;
  wire[3:0] T208;
  wire[7:0] T209;
  wire[3:0] T210;
  wire[3:0] T211;
  wire[15:0] T212;
  wire[7:0] T213;
  wire[3:0] T214;
  wire[3:0] T215;
  wire[7:0] T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[286:0] T453;
  wire[127:0] T219;
  wire[127:0] T220;
  wire[127:0] refill_data_0;
  wire[127:0] T221;
  wire[511:0] T222;
  wire[511:0] T223;
  wire[255:0] T224;
  reg [127:0] mem_tag_data_read_0;
  wire[127:0] T225;
  wire T226;
  wire T227;
  wire[3:0] T228;
  wire[1:0] T229;
  wire T230;
  reg [127:0] mem_tag_data_read_1;
  wire[127:0] T231;
  wire T232;
  wire T233;
  wire[255:0] T234;
  reg [127:0] mem_tag_data_read_2;
  wire[127:0] T235;
  wire T236;
  wire T237;
  reg [127:0] mem_tag_data_read_3;
  wire[127:0] T238;
  wire T239;
  wire T240;
  wire[127:0] refill_data_1;
  wire[127:0] T241;
  wire T242;
  wire[1:0] T243;
  wire[127:0] T244;
  wire[127:0] refill_data_2;
  wire[127:0] T245;
  wire[127:0] refill_data_3;
  wire[127:0] T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire[7:0] T253;
  wire[7:0] T254;
  wire[7:0] T255;
  wire[5:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire[5:0] T262;
  wire[16:0] T263;
  wire[15:0] T264;
  wire T265;
  wire[5:0] T266;
  wire[16:0] T267;
  wire[15:0] T268;
  wire T269;
  wire[127:0] T270;
  wire[127:0] T271;
  wire[127:0] T272;
  wire[127:0] mem_acq_data_write_0;
  wire[127:0] T273;
  wire[511:0] T274;
  wire[511:0] T275;
  wire[255:0] T276;
  wire[127:0] acq_data_no_tag_0;
  wire[127:0] T277;
  wire[63:0] T278;
  wire[63:0] T279;
  wire[127:0] acq_data_no_tag_1;
  wire[127:0] T280;
  wire[63:0] T281;
  wire[63:0] T282;
  wire[255:0] T283;
  wire[127:0] acq_data_no_tag_2;
  wire[127:0] T284;
  wire[63:0] T285;
  wire[63:0] T286;
  wire[127:0] acq_data_no_tag_3;
  wire[127:0] T287;
  wire[63:0] T288;
  wire[63:0] T289;
  wire[127:0] mem_acq_data_write_1;
  wire[127:0] T290;
  wire T291;
  wire[1:0] T292;
  wire[127:0] T293;
  wire[127:0] mem_acq_data_write_2;
  wire[127:0] T294;
  wire[127:0] mem_acq_data_write_3;
  wire[127:0] T295;
  wire T296;
  wire T297;
  wire[127:0] T298;
  wire[127:0] T299;
  wire[127:0] mem_tag_data_write_0;
  wire[127:0] T300;
  wire[511:0] T301;
  wire[511:0] T302;
  wire[255:0] T303;
  reg [127:0] wb_data_0;
  wire[127:0] T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[1:0] T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  reg [127:0] wb_data_1;
  wire[127:0] T313;
  wire T314;
  wire T315;
  wire[255:0] T316;
  reg [127:0] wb_data_2;
  wire[127:0] T317;
  wire T318;
  wire T319;
  reg [127:0] wb_data_3;
  wire[127:0] T320;
  wire T321;
  wire T322;
  wire[127:0] mem_tag_data_write_1;
  wire[127:0] T323;
  wire T324;
  wire[1:0] T325;
  wire[127:0] T326;
  wire[127:0] mem_tag_data_write_2;
  wire[127:0] T327;
  wire[127:0] mem_tag_data_write_3;
  wire[127:0] T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire[4:0] T454;
  wire[1:0] T338;
  wire[1:0] T339;
  wire[25:0] T340;
  wire[25:0] T341;
  wire[25:0] T342;
  wire[31:0] T343;
  wire[23:0] T344;
  wire[27:0] T345;
  wire[31:0] T346;
  wire[25:0] T347;
  wire[9:0] T348;
  wire[15:0] T349;
  reg [16:0] acq_repl_meta;
  wire[16:0] T350;
  wire[25:0] T351;
  wire[31:0] T352;
  wire[23:0] T353;
  wire[27:0] T354;
  wire[31:0] T355;
  wire T356;
  wire T357;
  wire[1:0] T358;
  wire T359;
  wire T360;
  wire[4:0] T361;
  reg [4:0] acq_src;
  wire[4:0] T362;
  wire[135:0] T363;
  wire[135:0] T364;
  wire[135:0] T365;
  wire[135:0] gnt_data_0;
  wire[135:0] T366;
  wire[543:0] T367;
  wire[543:0] T368;
  wire[271:0] T369;
  wire[135:0] T370;
  wire[67:0] T371;
  wire[63:0] T372;
  wire[511:0] T373;
  wire[511:0] T374;
  wire[255:0] T375;
  reg [127:0] mem_acq_data_read_0;
  wire[127:0] T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[1:0] T380;
  wire T381;
  reg [127:0] mem_acq_data_read_1;
  wire[127:0] T382;
  wire T383;
  wire T384;
  wire[255:0] T385;
  reg [127:0] mem_acq_data_read_2;
  wire[127:0] T386;
  wire T387;
  wire T388;
  reg [127:0] mem_acq_data_read_3;
  wire[127:0] T389;
  wire T390;
  wire T391;
  wire[3:0] T392;
  reg [31:0] gnt_tag;
  wire[31:0] T455;
  wire[127:0] T393;
  wire[127:0] T456;
  wire[127:0] T394;
  wire[7:0] T395;
  wire[1:0] T396;
  wire T397;
  wire[67:0] T398;
  wire[63:0] T399;
  wire[3:0] T400;
  wire[135:0] T401;
  wire[67:0] T402;
  wire[63:0] T403;
  wire[3:0] T404;
  wire[67:0] T405;
  wire[63:0] T406;
  wire[3:0] T407;
  wire[271:0] T408;
  wire[135:0] T409;
  wire[67:0] T410;
  wire[63:0] T411;
  wire[3:0] T412;
  wire[67:0] T413;
  wire[63:0] T414;
  wire[3:0] T415;
  wire[135:0] T416;
  wire[67:0] T417;
  wire[63:0] T418;
  wire[3:0] T419;
  wire[67:0] T420;
  wire[63:0] T421;
  wire[3:0] T422;
  wire[135:0] gnt_data_1;
  wire[135:0] T423;
  wire T424;
  wire[1:0] T425;
  wire[135:0] T426;
  wire[135:0] gnt_data_2;
  wire[135:0] T427;
  wire[135:0] gnt_data_3;
  wire[135:0] T428;
  wire T429;
  wire T430;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    collect_acq_data = {1{$random}};
    acq_data_cnt = {1{$random}};
    state = {1{$random}};
    acq_wr = {1{$random}};
    wb_read_cnt = {1{$random}};
    wb_data_cnt = {1{$random}};
    mem_tag_cmd_sent = {1{$random}};
    acq_data_process = {1{$random}};
    mem_acq_data_sent = {1{$random}};
    mem_acq_data_write_cnt = {1{$random}};
    mem_acq_cmd_sent = {1{$random}};
    mem_tag_data_sent = {1{$random}};
    mem_tag_data_write_cnt = {1{$random}};
    refill_data_cnt = {1{$random}};
    gnt_enable = {1{$random}};
    gnt_data_cnt = {1{$random}};
    mem_acq_gnt_ready = {1{$random}};
    mem_acq_data_read_cnt = {1{$random}};
    acq_addr = {1{$random}};
    mem_tag_refill_ready = {1{$random}};
    mem_tag_data_read_cnt = {1{$random}};
    acq_way_en = {1{$random}};
    acq_data_0 = {5{$random}};
    acq_data_1 = {5{$random}};
    acq_data_2 = {5{$random}};
    acq_data_3 = {5{$random}};
    mem_tag_data_read_0 = {4{$random}};
    mem_tag_data_read_1 = {4{$random}};
    mem_tag_data_read_2 = {4{$random}};
    mem_tag_data_read_3 = {4{$random}};
    wb_data_0 = {4{$random}};
    wb_data_1 = {4{$random}};
    wb_data_2 = {4{$random}};
    wb_data_3 = {4{$random}};
    acq_repl_meta = {1{$random}};
    acq_src = {1{$random}};
    mem_acq_data_read_0 = {4{$random}};
    mem_acq_data_read_1 = {4{$random}};
    mem_acq_data_read_2 = {4{$random}};
    mem_acq_data_read_3 = {4{$random}};
    gnt_tag = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_acq_match = T0;
  assign T0 = T149 & collect_acq_data;
  assign T431 = reset ? 1'h0 : T1;
  assign T1 = T147 ? acq_has_data : T2;
  assign T2 = T3 ? 1'h0 : collect_acq_data;
  assign T3 = T12 & acq_data_done;
  assign acq_data_done = T7 & T4;
  assign T4 = acq_data_cnt == 2'h3;
  assign T432 = reset ? 2'h0 : T5;
  assign T5 = T7 ? T6 : acq_data_cnt;
  assign T6 = acq_data_cnt + 2'h1;
  assign T7 = T11 & acq_has_data;
  assign T11 = io_uncached_acquire_ready & io_uncached_acquire_valid;
  assign T12 = collect_acq_data | T13;
  assign T13 = state == 4'h0;
  assign T433 = reset ? 4'h0 : T14;
  assign T14 = T123 ? 4'h0 : T15;
  assign T15 = T122 ? 4'he : T16;
  assign T16 = T120 ? T119 : T17;
  assign T17 = T111 ? 4'hc : T18;
  assign T18 = T107 ? 4'hb : T19;
  assign T19 = T62 ? 4'ha : T20;
  assign T20 = T55 ? 4'h9 : T21;
  assign T21 = T47 ? 4'h8 : T22;
  assign T22 = T45 ? 4'h7 : T23;
  assign T23 = T41 ? 4'he : T24;
  assign T24 = T40 ? 4'hd : T25;
  assign T25 = T38 ? 4'h4 : T26;
  assign T26 = T36 ? T31 : T27;
  assign T27 = T29 ? 4'h2 : T28;
  assign T28 = T147 ? 4'h1 : state;
  assign T29 = T30 & io_meta_read_ready;
  assign T30 = 4'h1 == state;
  assign T31 = io_meta_resp_bits_hit ? T34 : T32;
  assign T32 = T33 ? 4'h6 : 4'ha;
  assign T33 = io_meta_resp_bits_tag[5'h10:5'h10];
  assign T34 = acq_wr ? 4'h5 : 4'h3;
  assign T434 = reset ? 1'h0 : T35;
  assign T35 = T147 ? acq_has_data : acq_wr;
  assign T36 = T37 & io_meta_resp_valid;
  assign T37 = 4'h2 == state;
  assign T38 = T39 & io_data_read_ready;
  assign T39 = 4'h3 == state;
  assign T40 = 4'h4 == state;
  assign T41 = T42 & io_data_write_ready;
  assign T42 = T44 & T43;
  assign T43 = collect_acq_data ^ 1'h1;
  assign T44 = 4'h5 == state;
  assign T45 = T46 & io_data_read_ready;
  assign T46 = 4'h6 == state;
  assign T47 = T54 & wb_read_done;
  assign wb_read_done = T51 & T48;
  assign T48 = wb_read_cnt == 2'h3;
  assign T435 = reset ? 2'h0 : T49;
  assign T49 = T51 ? T50 : wb_read_cnt;
  assign T50 = wb_read_cnt + 2'h1;
  assign T51 = T53 & T52;
  assign T52 = state != 4'h3;
  assign T53 = io_data_read_ready & io_data_read_valid;
  assign T54 = 4'h7 == state;
  assign T55 = T61 & wb_data_done;
  assign wb_data_done = T59 & T56;
  assign T56 = wb_data_cnt == 2'h3;
  assign T436 = reset ? 2'h0 : T57;
  assign T57 = T59 ? T58 : wb_data_cnt;
  assign T58 = wb_data_cnt + 2'h1;
  assign T59 = io_data_resp_valid & T60;
  assign T60 = state != 4'h4;
  assign T61 = 4'h8 == state;
  assign T62 = T106 & T63;
  assign T63 = mem_tag_data_sent & mem_tag_cmd_sent;
  assign T437 = reset ? 1'h0 : T64;
  assign T64 = T62 ? 1'h0 : T65;
  assign T65 = T66 ? 1'h1 : mem_tag_cmd_sent;
  assign T66 = T67 & io_mem_req_cmd_ready;
  assign T67 = T69 & T68;
  assign T68 = mem_tag_cmd_sent ^ 1'h1;
  assign T69 = T94 & T70;
  assign T70 = acq_data_process ^ 1'h1;
  assign T438 = reset ? 1'h0 : T71;
  assign T71 = T147 ? 1'h1 : T72;
  assign T72 = T73 ? 1'h0 : acq_data_process;
  assign T73 = T92 & T74;
  assign T74 = mem_acq_cmd_sent & mem_acq_data_sent;
  assign T439 = reset ? 1'h0 : T75;
  assign T75 = T73 ? 1'h0 : T76;
  assign T76 = T77 ? 1'h1 : mem_acq_data_sent;
  assign T77 = T85 & T78;
  assign T78 = T84 | mem_acq_data_write_done;
  assign mem_acq_data_write_done = T82 & T79;
  assign T79 = mem_acq_data_write_cnt == 2'h3;
  assign T440 = reset ? 2'h0 : T80;
  assign T80 = T82 ? T81 : mem_acq_data_write_cnt;
  assign T81 = mem_acq_data_write_cnt + 2'h1;
  assign T82 = T83 & acq_data_process;
  assign T83 = io_mem_req_data_ready & io_mem_req_data_valid;
  assign T84 = acq_wr ^ 1'h1;
  assign T85 = T92 & T86;
  assign T86 = mem_acq_data_sent ^ 1'h1;
  assign T441 = reset ? 1'h0 : T87;
  assign T87 = T73 ? 1'h0 : T88;
  assign T88 = T89 ? 1'h1 : mem_acq_cmd_sent;
  assign T89 = T90 & io_mem_req_cmd_ready;
  assign T90 = T92 & T91;
  assign T91 = mem_acq_cmd_sent ^ 1'h1;
  assign T92 = acq_data_process & T93;
  assign T93 = collect_acq_data ^ 1'h1;
  assign T94 = state == 4'h9;
  assign T442 = reset ? 1'h0 : T95;
  assign T95 = T62 ? 1'h0 : T96;
  assign T96 = T97 ? 1'h1 : mem_tag_data_sent;
  assign T97 = T104 & mem_tag_data_write_done;
  assign mem_tag_data_write_done = T101 & T98;
  assign T98 = mem_tag_data_write_cnt == 2'h3;
  assign T443 = reset ? 2'h0 : T99;
  assign T99 = T101 ? T100 : mem_tag_data_write_cnt;
  assign T100 = mem_tag_data_write_cnt + 2'h1;
  assign T101 = T103 & T102;
  assign T102 = acq_data_process ^ 1'h1;
  assign T103 = io_mem_req_data_ready & io_mem_req_data_valid;
  assign T104 = T69 & T105;
  assign T105 = mem_tag_data_sent ^ 1'h1;
  assign T106 = 4'h9 == state;
  assign T107 = T108 & io_mem_req_cmd_ready;
  assign T108 = T110 & T109;
  assign T109 = acq_data_process ^ 1'h1;
  assign T110 = 4'ha == state;
  assign T111 = T118 & refill_data_done;
  assign refill_data_done = T115 & T112;
  assign T112 = refill_data_cnt == 2'h3;
  assign T444 = reset ? 2'h0 : T113;
  assign T113 = T115 ? T114 : refill_data_cnt;
  assign T114 = refill_data_cnt + 2'h1;
  assign T115 = T117 & T116;
  assign T116 = state == 4'hb;
  assign T117 = io_data_write_ready & io_data_write_valid;
  assign T118 = 4'hb == state;
  assign T119 = acq_wr ? 4'h5 : 4'h3;
  assign T120 = T121 & io_meta_write_ready;
  assign T121 = 4'hc == state;
  assign T122 = 4'hd == state;
  assign T123 = T146 & T124;
  assign T124 = T126 & T125;
  assign T125 = acq_data_process ^ 1'h1;
  assign T126 = gnt_enable ^ 1'h1;
  assign T445 = reset ? 1'h0 : T127;
  assign T127 = T122 ? 1'h1 : T128;
  assign T128 = T129 ? 1'h0 : gnt_enable;
  assign T129 = T136 & gnt_data_done;
  assign gnt_data_done = T133 & T130;
  assign T130 = gnt_data_cnt == 2'h3;
  assign T446 = reset ? 2'h0 : T131;
  assign T131 = T133 ? T132 : gnt_data_cnt;
  assign T132 = gnt_data_cnt + 2'h1;
  assign T133 = T135 & T134;
  assign T134 = acq_wr ^ 1'h1;
  assign T135 = io_uncached_grant_ready & io_uncached_grant_valid;
  assign T136 = gnt_enable & mem_acq_gnt_ready;
  assign T447 = reset ? 1'h0 : T137;
  assign T137 = T139 ? 1'h1 : T138;
  assign T138 = T129 ? 1'h0 : mem_acq_gnt_ready;
  assign T139 = io_mem_resp_valid & mem_acq_data_read_done;
  assign mem_acq_data_read_done = T143 & T140;
  assign T140 = mem_acq_data_read_cnt == 2'h3;
  assign T448 = reset ? 2'h0 : T141;
  assign T141 = T143 ? T142 : mem_acq_data_read_cnt;
  assign T142 = mem_acq_data_read_cnt + 2'h1;
  assign T143 = io_mem_resp_valid & mem_resp_is_acq;
  assign mem_resp_is_acq = T144;
  assign T144 = T145 == 1'h0;
  assign T145 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign T146 = 4'he == state;
  assign acq_has_data = io_uncached_acquire_bits_payload_uncached ? T8 : 1'h0;
  assign T8 = T10 | T9;
  assign T9 = 2'h2 == io_uncached_acquire_bits_payload_a_type;
  assign T10 = 2'h1 == io_uncached_acquire_bits_payload_a_type;
  assign T147 = T148 & io_uncached_acquire_valid;
  assign T148 = 4'h0 == state;
  assign T149 = acq_wr & T150;
  assign T150 = acq_addr == io_uncached_acquire_bits_payload_addr;
  assign T151 = T147 ? io_uncached_acquire_bits_payload_addr : acq_addr;
  assign io_acq_conflict = T152;
  assign T152 = T154 & T153;
  assign T153 = collect_acq_data ^ 1'h1;
  assign T154 = T156 & T155;
  assign T155 = state != 4'h0;
  assign T156 = T158 == T157;
  assign T157 = io_uncached_acquire_bits_payload_addr[4'h9:3'h4];
  assign T158 = acq_addr[4'h9:3'h4];
  assign io_data_write_bits_wmask = T159;
  assign T159 = T162 ? 4'hf : T160;
  assign T160 = 1'h1 << T161;
  assign T161 = acq_addr[1'h1:1'h0];
  assign T162 = T172 & mem_tag_refill_ready;
  assign T449 = reset ? 1'h0 : T163;
  assign T163 = T111 ? 1'h0 : T164;
  assign T164 = T165 ? 1'h1 : mem_tag_refill_ready;
  assign T165 = io_mem_resp_valid & mem_tag_data_read_done;
  assign mem_tag_data_read_done = T169 & T166;
  assign T166 = mem_tag_data_read_cnt == 2'h3;
  assign T450 = reset ? 2'h0 : T167;
  assign T167 = T169 ? T168 : mem_tag_data_read_cnt;
  assign T168 = mem_tag_data_read_cnt + 2'h1;
  assign T169 = io_mem_resp_valid & mem_resp_is_tag;
  assign mem_resp_is_tag = T170;
  assign T170 = T171 == 1'h1;
  assign T171 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign T172 = state == 4'hb;
  assign io_data_write_bits_way_en = acq_way_en;
  assign T451 = reset ? 8'h0 : T173;
  assign T173 = T174 ? io_meta_resp_bits_way_en : acq_way_en;
  assign T174 = T175 & io_meta_resp_valid;
  assign T175 = state == 4'h2;
  assign io_data_write_bits_addr = T176;
  assign T176 = T162 ? T178 : T177;
  assign T177 = acq_addr[4'h9:2'h2];
  assign T178 = {T179, refill_data_cnt};
  assign T179 = acq_addr[4'h9:3'h4];
  assign io_data_write_bits_data = T452;
  assign T452 = T180[7'h7f:1'h0];
  assign T180 = T162 ? T453 : T181;
  assign T181 = T184 << T182;
  assign T182 = T183 * 6'h20;
  assign T183 = acq_addr[1'h1:1'h0];
  assign T184 = T185;
  assign T185 = {T212, T186};
  assign T186 = {T209, T187};
  assign T187 = {T208, T188};
  assign T188 = T189[7'h43:7'h40];
  assign T189 = T190;
  assign T190 = {T201, T191};
  assign T191 = {acq_data_1, acq_data_0};
  assign T192 = T193 ? io_uncached_acquire_bits_payload_data : acq_data_0;
  assign T193 = T197 & T194;
  assign T194 = T195[1'h0:1'h0];
  assign T195 = 1'h1 << T196;
  assign T196 = acq_data_cnt;
  assign T197 = T12 & io_uncached_acquire_valid;
  assign T198 = T199 ? io_uncached_acquire_bits_payload_data : acq_data_1;
  assign T199 = T197 & T200;
  assign T200 = T195[1'h1:1'h1];
  assign T201 = {acq_data_3, acq_data_2};
  assign T202 = T203 ? io_uncached_acquire_bits_payload_data : acq_data_2;
  assign T203 = T197 & T204;
  assign T204 = T195[2'h2:2'h2];
  assign T205 = T206 ? io_uncached_acquire_bits_payload_data : acq_data_3;
  assign T206 = T197 & T207;
  assign T207 = T195[2'h3:2'h3];
  assign T208 = T189[8'h87:8'h84];
  assign T209 = {T211, T210};
  assign T210 = T189[8'hcb:8'hc8];
  assign T211 = T189[9'h10f:9'h10c];
  assign T212 = {T216, T213};
  assign T213 = {T215, T214};
  assign T214 = T189[9'h153:9'h150];
  assign T215 = T189[9'h197:9'h194];
  assign T216 = {T218, T217};
  assign T217 = T189[9'h1db:9'h1d8];
  assign T218 = T189[10'h21f:10'h21c];
  assign T453 = {159'h0, T219};
  assign T219 = T248 ? T244 : T220;
  assign T220 = T242 ? refill_data_1 : refill_data_0;
  assign refill_data_0 = T221;
  assign T221 = T222[7'h7f:1'h0];
  assign T222 = T223;
  assign T223 = {T234, T224};
  assign T224 = {mem_tag_data_read_1, mem_tag_data_read_0};
  assign T225 = T226 ? io_mem_resp_bits_data : mem_tag_data_read_0;
  assign T226 = T230 & T227;
  assign T227 = T228[1'h0:1'h0];
  assign T228 = 1'h1 << T229;
  assign T229 = mem_tag_data_read_cnt;
  assign T230 = io_mem_resp_valid & mem_resp_is_tag;
  assign T231 = T232 ? io_mem_resp_bits_data : mem_tag_data_read_1;
  assign T232 = T230 & T233;
  assign T233 = T228[1'h1:1'h1];
  assign T234 = {mem_tag_data_read_3, mem_tag_data_read_2};
  assign T235 = T236 ? io_mem_resp_bits_data : mem_tag_data_read_2;
  assign T236 = T230 & T237;
  assign T237 = T228[2'h2:2'h2];
  assign T238 = T239 ? io_mem_resp_bits_data : mem_tag_data_read_3;
  assign T239 = T230 & T240;
  assign T240 = T228[2'h3:2'h3];
  assign refill_data_1 = T241;
  assign T241 = T222[8'hff:8'h80];
  assign T242 = T243[1'h0:1'h0];
  assign T243 = refill_data_cnt;
  assign T244 = T247 ? refill_data_3 : refill_data_2;
  assign refill_data_2 = T245;
  assign T245 = T222[9'h17f:9'h100];
  assign refill_data_3 = T246;
  assign T246 = T222[9'h1ff:9'h180];
  assign T247 = T243[1'h0:1'h0];
  assign T248 = T243[1'h1:1'h1];
  assign io_data_write_valid = T249;
  assign T249 = T162 ? 1'h1 : T250;
  assign T250 = T252 & T251;
  assign T251 = collect_acq_data ^ 1'h1;
  assign T252 = state == 4'h5;
  assign io_data_read_bits_way_en = acq_way_en;
  assign io_data_read_bits_addr = T253;
  assign T253 = T257 ? T255 : T254;
  assign T254 = acq_addr[4'h9:2'h2];
  assign T255 = {T256, wb_read_cnt};
  assign T256 = acq_addr[4'h9:3'h4];
  assign T257 = T259 | T258;
  assign T258 = state == 4'h7;
  assign T259 = state == 4'h6;
  assign io_data_read_bits_id = 1'h0;
  assign io_data_read_valid = T260;
  assign T260 = T257 ? 1'h1 : T261;
  assign T261 = state == 4'h3;
  assign io_meta_write_bits_way_en = acq_way_en;
  assign io_meta_write_bits_idx = T262;
  assign T262 = acq_addr[4'h9:3'h4];
  assign io_meta_write_bits_tag = T263;
  assign T263 = {1'h1, T264};
  assign T264 = acq_addr >> 4'ha;
  assign io_meta_write_valid = T265;
  assign T265 = state == 4'hc;
  assign io_meta_read_bits_idx = T266;
  assign T266 = acq_addr[4'h9:3'h4];
  assign io_meta_read_bits_tag = T267;
  assign T267 = {1'h1, T268};
  assign T268 = acq_addr >> 4'ha;
  assign io_meta_read_bits_id = 1'h0;
  assign io_meta_read_valid = T269;
  assign T269 = state == 4'h1;
  assign io_mem_req_data_bits_data = T270;
  assign T270 = T104 ? T298 : T271;
  assign T271 = T297 ? T293 : T272;
  assign T272 = T291 ? mem_acq_data_write_1 : mem_acq_data_write_0;
  assign mem_acq_data_write_0 = T273;
  assign T273 = T274[7'h7f:1'h0];
  assign T274 = T275;
  assign T275 = {T283, T276};
  assign T276 = {acq_data_no_tag_1, acq_data_no_tag_0};
  assign acq_data_no_tag_0 = T277;
  assign T277 = {T279, T278};
  assign T278 = acq_data_0[6'h3f:1'h0];
  assign T279 = acq_data_0[8'h83:7'h44];
  assign acq_data_no_tag_1 = T280;
  assign T280 = {T282, T281};
  assign T281 = acq_data_1[6'h3f:1'h0];
  assign T282 = acq_data_1[8'h83:7'h44];
  assign T283 = {acq_data_no_tag_3, acq_data_no_tag_2};
  assign acq_data_no_tag_2 = T284;
  assign T284 = {T286, T285};
  assign T285 = acq_data_2[6'h3f:1'h0];
  assign T286 = acq_data_2[8'h83:7'h44];
  assign acq_data_no_tag_3 = T287;
  assign T287 = {T289, T288};
  assign T288 = acq_data_3[6'h3f:1'h0];
  assign T289 = acq_data_3[8'h83:7'h44];
  assign mem_acq_data_write_1 = T290;
  assign T290 = T274[8'hff:8'h80];
  assign T291 = T292[1'h0:1'h0];
  assign T292 = mem_acq_data_write_cnt;
  assign T293 = T296 ? mem_acq_data_write_3 : mem_acq_data_write_2;
  assign mem_acq_data_write_2 = T294;
  assign T294 = T274[9'h17f:9'h100];
  assign mem_acq_data_write_3 = T295;
  assign T295 = T274[9'h1ff:9'h180];
  assign T296 = T292[1'h0:1'h0];
  assign T297 = T292[1'h1:1'h1];
  assign T298 = T330 ? T326 : T299;
  assign T299 = T324 ? mem_tag_data_write_1 : mem_tag_data_write_0;
  assign mem_tag_data_write_0 = T300;
  assign T300 = T301[7'h7f:1'h0];
  assign T301 = T302;
  assign T302 = {T316, T303};
  assign T303 = {wb_data_1, wb_data_0};
  assign T304 = T305 ? io_data_resp_bits_data : wb_data_0;
  assign T305 = T309 & T306;
  assign T306 = T307[1'h0:1'h0];
  assign T307 = 1'h1 << T308;
  assign T308 = wb_data_cnt;
  assign T309 = T310 & io_data_resp_valid;
  assign T310 = T312 | T311;
  assign T311 = state == 4'h8;
  assign T312 = state == 4'h7;
  assign T313 = T314 ? io_data_resp_bits_data : wb_data_1;
  assign T314 = T309 & T315;
  assign T315 = T307[1'h1:1'h1];
  assign T316 = {wb_data_3, wb_data_2};
  assign T317 = T318 ? io_data_resp_bits_data : wb_data_2;
  assign T318 = T309 & T319;
  assign T319 = T307[2'h2:2'h2];
  assign T320 = T321 ? io_data_resp_bits_data : wb_data_3;
  assign T321 = T309 & T322;
  assign T322 = T307[2'h3:2'h3];
  assign mem_tag_data_write_1 = T323;
  assign T323 = T301[8'hff:8'h80];
  assign T324 = T325[1'h0:1'h0];
  assign T325 = mem_tag_data_write_cnt;
  assign T326 = T329 ? mem_tag_data_write_3 : mem_tag_data_write_2;
  assign mem_tag_data_write_2 = T327;
  assign T327 = T301[9'h17f:9'h100];
  assign mem_tag_data_write_3 = T328;
  assign T328 = T301[9'h1ff:9'h180];
  assign T329 = T325[1'h0:1'h0];
  assign T330 = T325[1'h1:1'h1];
  assign io_mem_req_data_valid = T331;
  assign T331 = T104 ? 1'h1 : T332;
  assign T332 = T85 & acq_wr;
  assign io_mem_req_cmd_bits_rw = T333;
  assign T333 = T335 ? 1'h0 : T334;
  assign T334 = T67 ? 1'h1 : acq_wr;
  assign T335 = T337 & T336;
  assign T336 = acq_data_process ^ 1'h1;
  assign T337 = state == 4'ha;
  assign io_mem_req_cmd_bits_tag = T454;
  assign T454 = {3'h0, T338};
  assign T338 = T335 ? 2'h1 : T339;
  assign T339 = T67 ? 2'h1 : 2'h0;
  assign io_mem_req_cmd_bits_addr = T340;
  assign T340 = T335 ? T351 : T341;
  assign T341 = T67 ? T342 : acq_addr;
  assign T342 = T343 >> 3'h6;
  assign T343 = {8'hf, T344};
  assign T344 = T345[5'h17:1'h0];
  assign T345 = T346 >> 3'h4;
  assign T346 = {T347, 6'h0};
  assign T347 = {T349, T348};
  assign T348 = acq_addr[4'h9:1'h0];
  assign T349 = acq_repl_meta[4'hf:1'h0];
  assign T350 = T174 ? io_meta_resp_bits_tag : acq_repl_meta;
  assign T351 = T352 >> 3'h6;
  assign T352 = {8'hf, T353};
  assign T353 = T354[5'h17:1'h0];
  assign T354 = T355 >> 3'h4;
  assign T355 = {acq_addr, 6'h0};
  assign io_mem_req_cmd_valid = T356;
  assign T356 = T335 ? 1'h1 : T357;
  assign T357 = T67 ? 1'h1 : T90;
//  assign io_uncached_finish_ready = {1{$random}};
  assign io_uncached_grant_bits_payload_g_type = T358;
  assign T358 = 2'h0;
  assign io_uncached_grant_bits_payload_uncached = T359;
  assign T359 = 1'h1;
  assign io_uncached_grant_bits_payload_manager_xact_id = T360;
  assign T360 = 1'h0;
  assign io_uncached_grant_bits_payload_client_xact_id = T361;
  assign T361 = acq_src;
  assign T362 = T147 ? io_uncached_acquire_bits_payload_client_xact_id : acq_src;
  assign io_uncached_grant_bits_payload_data = T363;
  assign T363 = T364;
  assign T364 = T430 ? T426 : T365;
  assign T365 = T424 ? gnt_data_1 : gnt_data_0;
  assign gnt_data_0 = T366;
  assign T366 = T367[8'h87:1'h0];
  assign T367 = T368;
  assign T368 = {T408, T369};
  assign T369 = {T401, T370};
  assign T370 = {T398, T371};
  assign T371 = {T392, T372};
  assign T372 = T373[6'h3f:1'h0];
  assign T373 = T374;
  assign T374 = {T385, T375};
  assign T375 = {mem_acq_data_read_1, mem_acq_data_read_0};
  assign T376 = T377 ? io_mem_resp_bits_data : mem_acq_data_read_0;
  assign T377 = T381 & T378;
  assign T378 = T379[1'h0:1'h0];
  assign T379 = 1'h1 << T380;
  assign T380 = mem_acq_data_read_cnt;
  assign T381 = io_mem_resp_valid & mem_resp_is_acq;
  assign T382 = T383 ? io_mem_resp_bits_data : mem_acq_data_read_1;
  assign T383 = T381 & T384;
  assign T384 = T379[1'h1:1'h1];
  assign T385 = {mem_acq_data_read_3, mem_acq_data_read_2};
  assign T386 = T387 ? io_mem_resp_bits_data : mem_acq_data_read_2;
  assign T387 = T381 & T388;
  assign T388 = T379[2'h2:2'h2];
  assign T389 = T390 ? io_mem_resp_bits_data : mem_acq_data_read_3;
  assign T390 = T381 & T391;
  assign T391 = T379[2'h3:2'h3];
  assign T392 = gnt_tag[2'h3:1'h0];
  assign T455 = T393[5'h1f:1'h0];
  assign T393 = T397 ? T394 : T456;
  assign T456 = {96'h0, gnt_tag};
  assign T394 = io_data_resp_bits_data >> T395;
  assign T395 = T396 * 6'h20;
  assign T396 = acq_addr[1'h1:1'h0];
  assign T397 = state == 4'h4;
  assign T398 = {T400, T399};
  assign T399 = T373[7'h7f:7'h40];
  assign T400 = gnt_tag[3'h7:3'h4];
  assign T401 = {T405, T402};
  assign T402 = {T404, T403};
  assign T403 = T373[8'hbf:8'h80];
  assign T404 = gnt_tag[4'hb:4'h8];
  assign T405 = {T407, T406};
  assign T406 = T373[8'hff:8'hc0];
  assign T407 = gnt_tag[4'hf:4'hc];
  assign T408 = {T416, T409};
  assign T409 = {T413, T410};
  assign T410 = {T412, T411};
  assign T411 = T373[9'h13f:9'h100];
  assign T412 = gnt_tag[5'h13:5'h10];
  assign T413 = {T415, T414};
  assign T414 = T373[9'h17f:9'h140];
  assign T415 = gnt_tag[5'h17:5'h14];
  assign T416 = {T420, T417};
  assign T417 = {T419, T418};
  assign T418 = T373[9'h1bf:9'h180];
  assign T419 = gnt_tag[5'h1b:5'h18];
  assign T420 = {T422, T421};
  assign T421 = T373[9'h1ff:9'h1c0];
  assign T422 = gnt_tag[5'h1f:5'h1c];
  assign gnt_data_1 = T423;
  assign T423 = T367[9'h10f:8'h88];
  assign T424 = T425[1'h0:1'h0];
  assign T425 = gnt_data_cnt;
  assign T426 = T429 ? gnt_data_3 : gnt_data_2;
  assign gnt_data_2 = T427;
  assign T427 = T367[9'h197:9'h110];
  assign gnt_data_3 = T428;
  assign T428 = T367[10'h21f:9'h198];
  assign T429 = T425[1'h0:1'h0];
  assign T430 = T425[1'h1:1'h1];
//  assign io_uncached_grant_bits_header_dst = {1{$random}};
//  assign io_uncached_grant_bits_header_src = {1{$random}};
  assign io_uncached_grant_valid = T136;
  assign io_uncached_acquire_ready = T12;

  always @(posedge clk) begin
    if(reset) begin
      collect_acq_data <= 1'h0;
    end else if(T147) begin
      collect_acq_data <= acq_has_data;
    end else if(T3) begin
      collect_acq_data <= 1'h0;
    end
    if(reset) begin
      acq_data_cnt <= 2'h0;
    end else if(T7) begin
      acq_data_cnt <= T6;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T123) begin
      state <= 4'h0;
    end else if(T122) begin
      state <= 4'he;
    end else if(T120) begin
      state <= T119;
    end else if(T111) begin
      state <= 4'hc;
    end else if(T107) begin
      state <= 4'hb;
    end else if(T62) begin
      state <= 4'ha;
    end else if(T55) begin
      state <= 4'h9;
    end else if(T47) begin
      state <= 4'h8;
    end else if(T45) begin
      state <= 4'h7;
    end else if(T41) begin
      state <= 4'he;
    end else if(T40) begin
      state <= 4'hd;
    end else if(T38) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= T31;
    end else if(T29) begin
      state <= 4'h2;
    end else if(T147) begin
      state <= 4'h1;
    end
    if(reset) begin
      acq_wr <= 1'h0;
    end else if(T147) begin
      acq_wr <= acq_has_data;
    end
    if(reset) begin
      wb_read_cnt <= 2'h0;
    end else if(T51) begin
      wb_read_cnt <= T50;
    end
    if(reset) begin
      wb_data_cnt <= 2'h0;
    end else if(T59) begin
      wb_data_cnt <= T58;
    end
    if(reset) begin
      mem_tag_cmd_sent <= 1'h0;
    end else if(T62) begin
      mem_tag_cmd_sent <= 1'h0;
    end else if(T66) begin
      mem_tag_cmd_sent <= 1'h1;
    end
    if(reset) begin
      acq_data_process <= 1'h0;
    end else if(T147) begin
      acq_data_process <= 1'h1;
    end else if(T73) begin
      acq_data_process <= 1'h0;
    end
    if(reset) begin
      mem_acq_data_sent <= 1'h0;
    end else if(T73) begin
      mem_acq_data_sent <= 1'h0;
    end else if(T77) begin
      mem_acq_data_sent <= 1'h1;
    end
    if(reset) begin
      mem_acq_data_write_cnt <= 2'h0;
    end else if(T82) begin
      mem_acq_data_write_cnt <= T81;
    end
    if(reset) begin
      mem_acq_cmd_sent <= 1'h0;
    end else if(T73) begin
      mem_acq_cmd_sent <= 1'h0;
    end else if(T89) begin
      mem_acq_cmd_sent <= 1'h1;
    end
    if(reset) begin
      mem_tag_data_sent <= 1'h0;
    end else if(T62) begin
      mem_tag_data_sent <= 1'h0;
    end else if(T97) begin
      mem_tag_data_sent <= 1'h1;
    end
    if(reset) begin
      mem_tag_data_write_cnt <= 2'h0;
    end else if(T101) begin
      mem_tag_data_write_cnt <= T100;
    end
    if(reset) begin
      refill_data_cnt <= 2'h0;
    end else if(T115) begin
      refill_data_cnt <= T114;
    end
    if(reset) begin
      gnt_enable <= 1'h0;
    end else if(T122) begin
      gnt_enable <= 1'h1;
    end else if(T129) begin
      gnt_enable <= 1'h0;
    end
    if(reset) begin
      gnt_data_cnt <= 2'h0;
    end else if(T133) begin
      gnt_data_cnt <= T132;
    end
    if(reset) begin
      mem_acq_gnt_ready <= 1'h0;
    end else if(T139) begin
      mem_acq_gnt_ready <= 1'h1;
    end else if(T129) begin
      mem_acq_gnt_ready <= 1'h0;
    end
    if(reset) begin
      mem_acq_data_read_cnt <= 2'h0;
    end else if(T143) begin
      mem_acq_data_read_cnt <= T142;
    end
    if(T147) begin
      acq_addr <= io_uncached_acquire_bits_payload_addr;
    end
    if(reset) begin
      mem_tag_refill_ready <= 1'h0;
    end else if(T111) begin
      mem_tag_refill_ready <= 1'h0;
    end else if(T165) begin
      mem_tag_refill_ready <= 1'h1;
    end
    if(reset) begin
      mem_tag_data_read_cnt <= 2'h0;
    end else if(T169) begin
      mem_tag_data_read_cnt <= T168;
    end
    if(reset) begin
      acq_way_en <= 8'h0;
    end else if(T174) begin
      acq_way_en <= io_meta_resp_bits_way_en;
    end
    if(T193) begin
      acq_data_0 <= io_uncached_acquire_bits_payload_data;
    end
    if(T199) begin
      acq_data_1 <= io_uncached_acquire_bits_payload_data;
    end
    if(T203) begin
      acq_data_2 <= io_uncached_acquire_bits_payload_data;
    end
    if(T206) begin
      acq_data_3 <= io_uncached_acquire_bits_payload_data;
    end
    if(T226) begin
      mem_tag_data_read_0 <= io_mem_resp_bits_data;
    end
    if(T232) begin
      mem_tag_data_read_1 <= io_mem_resp_bits_data;
    end
    if(T236) begin
      mem_tag_data_read_2 <= io_mem_resp_bits_data;
    end
    if(T239) begin
      mem_tag_data_read_3 <= io_mem_resp_bits_data;
    end
    if(T305) begin
      wb_data_0 <= io_data_resp_bits_data;
    end
    if(T314) begin
      wb_data_1 <= io_data_resp_bits_data;
    end
    if(T318) begin
      wb_data_2 <= io_data_resp_bits_data;
    end
    if(T321) begin
      wb_data_3 <= io_data_resp_bits_data;
    end
    if(T174) begin
      acq_repl_meta <= io_meta_resp_bits_tag;
    end
    if(T147) begin
      acq_src <= io_uncached_acquire_bits_payload_client_xact_id;
    end
    if(T377) begin
      mem_acq_data_read_0 <= io_mem_resp_bits_data;
    end
    if(T383) begin
      mem_acq_data_read_1 <= io_mem_resp_bits_data;
    end
    if(T387) begin
      mem_acq_data_read_2 <= io_mem_resp_bits_data;
    end
    if(T390) begin
      mem_acq_data_read_3 <= io_mem_resp_bits_data;
    end
    gnt_tag <= T455;
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [4:0] io_enq_bits_payload_client_xact_id,
    input [135:0] io_enq_bits_payload_data,
    input  io_enq_bits_payload_uncached,
    input [1:0] io_enq_bits_payload_a_type,
    input [128:0] io_enq_bits_payload_subblock,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[4:0] io_deq_bits_payload_client_xact_id,
    output[135:0] io_deq_bits_payload_data,
    output io_deq_bits_payload_uncached,
    output[1:0] io_deq_bits_payload_a_type,
    output[128:0] io_deq_bits_payload_subblock,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T31;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T32;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[128:0] T10;
  wire[302:0] T11;
  reg [302:0] ram [7:0];
  wire[302:0] T12;
  wire[302:0] T13;
  wire[302:0] T14;
  wire[267:0] T15;
  wire[130:0] T16;
  wire[136:0] T17;
  wire[34:0] T18;
  wire[30:0] T19;
  wire[3:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[135:0] T23;
  wire[4:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {10{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_subblock = T10;
  assign T10 = T11[8'h80:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_a_type, io_enq_bits_payload_subblock};
  assign T17 = {io_enq_bits_payload_data, io_enq_bits_payload_uncached};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_a_type = T21;
  assign T21 = T11[8'h82:8'h81];
  assign io_deq_bits_payload_uncached = T22;
  assign T22 = T11[8'h83:8'h83];
  assign io_deq_bits_payload_data = T23;
  assign T23 = T11[9'h10b:8'h84];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T11[9'h110:9'h10c];
  assign io_deq_bits_payload_addr = T25;
  assign T25 = T11[9'h12a:9'h111];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[9'h12c:9'h12b];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[9'h12e:9'h12d];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T21;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T22;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  reg [31:0] ram [7:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[5:0] T15;
  wire[4:0] T16;
  wire[25:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_rw = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_addr, T15};
  assign T15 = {io_enq_bits_tag, io_enq_bits_rw};
  assign io_deq_bits_tag = T16;
  assign T16 = T11[3'h5:1'h1];
  assign io_deq_bits_addr = T17;
  assign T17 = T11[5'h1f:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T16;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T17;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T18;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[127:0] T11;
  reg [127:0] ram [7:0];
  wire[127:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T16 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T17 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T18 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_data;
  end
endmodule

module Arbiter_11(
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits = io_in_0_bits;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [135:0] io_in_0_bits_payload_data,
    input [4:0] io_in_0_bits_payload_client_xact_id,
    input  io_in_0_bits_payload_manager_xact_id,
    input  io_in_0_bits_payload_uncached,
    input [1:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[135:0] io_out_bits_payload_data,
    output[4:0] io_out_bits_payload_client_xact_id,
    output io_out_bits_payload_manager_xact_id,
    output io_out_bits_payload_uncached,
    output[1:0] io_out_bits_payload_g_type,
    output io_chosen
);

  wire chosen;
  wire T0;
  reg  lockIdx;
  wire T28;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg  locked;
  wire T29;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] T15;
  reg [1:0] R16;
  wire[1:0] T30;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  reg  last_grant;
  wire T31;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R16 = {1{$random}};
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : 1'h0;
  assign T28 = reset ? 1'h0 : T1;
  assign T1 = T2 ? 1'h0 : lockIdx;
  assign T2 = T4 & T3;
  assign T3 = locked ^ 1'h1;
  assign T4 = T10 & T5;
  assign T5 = io_out_bits_payload_uncached ? T7 : T6;
  assign T6 = 2'h1 == io_out_bits_payload_g_type;
  assign T7 = T9 | T8;
  assign T8 = 2'h2 == io_out_bits_payload_g_type;
  assign T9 = 2'h0 == io_out_bits_payload_g_type;
  assign T10 = io_out_ready & io_out_valid;
  assign T29 = reset ? 1'h0 : T11;
  assign T11 = T13 ? 1'h0 : T12;
  assign T12 = T2 ? 1'h1 : locked;
  assign T13 = T10 & T14;
  assign T14 = T15 == 2'h0;
  assign T15 = R16 + 2'h1;
  assign T30 = reset ? 2'h0 : T17;
  assign T17 = T4 ? T15 : R16;
  assign io_out_bits_payload_g_type = io_in_0_bits_payload_g_type;
  assign io_out_bits_payload_uncached = io_in_0_bits_payload_uncached;
  assign io_out_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign io_out_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_data = io_in_0_bits_payload_data;
  assign io_out_bits_header_dst = io_in_0_bits_header_dst;
  assign io_out_bits_header_src = io_in_0_bits_header_src;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T18;
  assign T18 = T19 & io_out_ready;
  assign T19 = locked ? T27 : T20;
  assign T20 = T26 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = io_in_0_valid & T23;
  assign T23 = last_grant < 1'h0;
  assign T31 = reset ? 1'h0 : T24;
  assign T24 = T25 ? chosen : last_grant;
  assign T25 = io_out_ready & io_out_valid;
  assign T26 = last_grant < 1'h0;
  assign T27 = lockIdx == 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h0;
    end else if(T2) begin
      lockIdx <= 1'h0;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T13) begin
      locked <= 1'h0;
    end else if(T2) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R16 <= 2'h0;
    end else if(T4) begin
      R16 <= T15;
    end
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T25) begin
      last_grant <= chosen;
    end
  end
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [4:0] io_in_0_bits_tag,
    input  io_in_0_bits_rw,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[4:0] io_out_bits_tag,
    output io_out_bits_rw,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  last_grant;
  wire T8;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_rw = io_in_0_bits_rw;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T0;
  assign T0 = T1 & io_out_ready;
  assign T1 = T7 | T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_0_valid & T4;
  assign T4 = last_grant < 1'h0;
  assign T8 = reset ? 1'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = last_grant < 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  reg  lockIdx;
  wire T22;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  locked;
  wire T23;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[1:0] T9;
  reg [1:0] R10;
  wire[1:0] T24;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  last_grant;
  wire T25;
  wire T18;
  wire T19;
  wire T20;
  wire T21;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R10 = {1{$random}};
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : 1'h0;
  assign T22 = reset ? 1'h0 : T1;
  assign T1 = T2 ? 1'h0 : lockIdx;
  assign T2 = T4 & T3;
  assign T3 = locked ^ 1'h1;
  assign T4 = io_out_ready & io_out_valid;
  assign T23 = reset ? 1'h0 : T5;
  assign T5 = T7 ? 1'h0 : T6;
  assign T6 = T2 ? 1'h1 : locked;
  assign T7 = T4 & T8;
  assign T8 = T9 == 2'h0;
  assign T9 = R10 + 2'h1;
  assign T24 = reset ? 2'h0 : T11;
  assign T11 = T4 ? T9 : R10;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = locked ? T21 : T14;
  assign T14 = T20 | T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T25 = reset ? 1'h0 : T18;
  assign T18 = T19 ? chosen : last_grant;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = last_grant < 1'h0;
  assign T21 = lockIdx == 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h0;
    end else if(T2) begin
      lockIdx <= 1'h0;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T7) begin
      locked <= 1'h0;
    end else if(T2) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R10 <= 2'h0;
    end else if(T4) begin
      R10 <= T9;
    end
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T19) begin
      last_grant <= chosen;
    end
  end
endmodule

module LockingRRArbiter_5(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_id,
    input [16:0] io_in_0_bits_tag,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_id,
    output[16:0] io_out_bits_tag,
    output[5:0] io_out_bits_idx,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  last_grant;
  wire T8;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_idx = io_in_0_bits_idx;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_id = io_in_0_bits_id;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T0;
  assign T0 = T1 & io_out_ready;
  assign T1 = T7 | T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_0_valid & T4;
  assign T4 = last_grant < 1'h0;
  assign T8 = reset ? 1'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = last_grant < 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module LockingRRArbiter_6(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [16:0] io_in_0_bits_tag,
    input [5:0] io_in_0_bits_idx,
    input [7:0] io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output[16:0] io_out_bits_tag,
    output[5:0] io_out_bits_idx,
    output[7:0] io_out_bits_way_en,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  last_grant;
  wire T8;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_way_en = io_in_0_bits_way_en;
  assign io_out_bits_idx = io_in_0_bits_idx;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T0;
  assign T0 = T1 & io_out_ready;
  assign T1 = T7 | T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_0_valid & T4;
  assign T4 = last_grant < 1'h0;
  assign T8 = reset ? 1'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = last_grant < 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module LockingRRArbiter_7(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_id,
    input [7:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_id,
    output[7:0] io_out_bits_addr,
    output[7:0] io_out_bits_way_en,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  last_grant;
  wire T8;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_way_en = io_in_0_bits_way_en;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_bits_id = io_in_0_bits_id;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T0;
  assign T0 = T1 & io_out_ready;
  assign T1 = T7 | T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_0_valid & T4;
  assign T4 = last_grant < 1'h0;
  assign T8 = reset ? 1'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = last_grant < 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module LockingRRArbiter_8(input clk, input reset,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [127:0] io_in_0_bits_data,
    input [7:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_way_en,
    input [3:0] io_in_0_bits_wmask,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[7:0] io_out_bits_addr,
    output[7:0] io_out_bits_way_en,
    output[3:0] io_out_bits_wmask,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  last_grant;
  wire T8;
  wire T5;
  wire T6;
  wire T7;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_wmask = io_in_0_bits_wmask;
  assign io_out_bits_way_en = io_in_0_bits_way_en;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = T0;
  assign T0 = T1 & io_out_ready;
  assign T1 = T7 | T2;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_in_0_valid & T4;
  assign T4 = last_grant < 1'h0;
  assign T8 = reset ? 1'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = last_grant < 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module TagCache(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [4:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [135:0] io_uncached_acquire_bits_payload_data,
    input  io_uncached_acquire_bits_payload_uncached,
    input [1:0] io_uncached_acquire_bits_payload_a_type,
    input [128:0] io_uncached_acquire_bits_payload_subblock,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    output[1:0] io_uncached_grant_bits_header_src,
    output[1:0] io_uncached_grant_bits_header_dst,
    output[135:0] io_uncached_grant_bits_payload_data,
    output[4:0] io_uncached_grant_bits_payload_client_xact_id,
    output io_uncached_grant_bits_payload_manager_xact_id,
    output io_uncached_grant_bits_payload_uncached,
    output[1:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input  io_uncached_finish_bits_payload_manager_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire T0;
  wire T1;
  wire acq_conflict;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire T12;
  wire T13;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire meta_io_resp_valid;
  wire meta_io_resp_bits_id;
  wire[16:0] meta_io_resp_bits_tag;
  wire meta_io_resp_bits_hit;
  wire[7:0] meta_io_resp_bits_way_en;
  wire data_io_read_ready;
  wire data_io_write_ready;
  wire data_io_resp_valid;
  wire data_io_resp_bits_id;
  wire[127:0] data_io_resp_bits_data;
  wire TagCacheTracker_io_uncached_acquire_ready;
  wire TagCacheTracker_io_uncached_grant_valid;
  wire[135:0] TagCacheTracker_io_uncached_grant_bits_payload_data;
  wire[4:0] TagCacheTracker_io_uncached_grant_bits_payload_client_xact_id;
  wire TagCacheTracker_io_uncached_grant_bits_payload_manager_xact_id;
  wire TagCacheTracker_io_uncached_grant_bits_payload_uncached;
  wire[1:0] TagCacheTracker_io_uncached_grant_bits_payload_g_type;
  wire TagCacheTracker_io_mem_req_cmd_valid;
  wire[25:0] TagCacheTracker_io_mem_req_cmd_bits_addr;
  wire[4:0] TagCacheTracker_io_mem_req_cmd_bits_tag;
  wire TagCacheTracker_io_mem_req_cmd_bits_rw;
  wire TagCacheTracker_io_mem_req_data_valid;
  wire[127:0] TagCacheTracker_io_mem_req_data_bits_data;
  wire TagCacheTracker_io_meta_read_valid;
  wire TagCacheTracker_io_meta_read_bits_id;
  wire[16:0] TagCacheTracker_io_meta_read_bits_tag;
  wire[5:0] TagCacheTracker_io_meta_read_bits_idx;
  wire TagCacheTracker_io_meta_write_valid;
  wire[16:0] TagCacheTracker_io_meta_write_bits_tag;
  wire[5:0] TagCacheTracker_io_meta_write_bits_idx;
  wire[7:0] TagCacheTracker_io_meta_write_bits_way_en;
  wire TagCacheTracker_io_data_read_valid;
  wire TagCacheTracker_io_data_read_bits_id;
  wire[7:0] TagCacheTracker_io_data_read_bits_addr;
  wire[7:0] TagCacheTracker_io_data_read_bits_way_en;
  wire TagCacheTracker_io_data_write_valid;
  wire[127:0] TagCacheTracker_io_data_write_bits_data;
  wire[7:0] TagCacheTracker_io_data_write_bits_addr;
  wire[7:0] TagCacheTracker_io_data_write_bits_way_en;
  wire[3:0] TagCacheTracker_io_data_write_bits_wmask;
  wire TagCacheTracker_io_acq_conflict;
  wire acqQueue_io_enq_ready;
  wire acqQueue_io_deq_valid;
  wire[1:0] acqQueue_io_deq_bits_header_src;
  wire[1:0] acqQueue_io_deq_bits_header_dst;
  wire[25:0] acqQueue_io_deq_bits_payload_addr;
  wire[4:0] acqQueue_io_deq_bits_payload_client_xact_id;
  wire[135:0] acqQueue_io_deq_bits_payload_data;
  wire acqQueue_io_deq_bits_payload_uncached;
  wire[1:0] acqQueue_io_deq_bits_payload_a_type;
  wire[128:0] acqQueue_io_deq_bits_payload_subblock;
  wire memCMDQueue_io_enq_ready;
  wire memCMDQueue_io_deq_valid;
  wire[25:0] memCMDQueue_io_deq_bits_addr;
  wire[4:0] memCMDQueue_io_deq_bits_tag;
  wire memCMDQueue_io_deq_bits_rw;
  wire memDataQueue_io_enq_ready;
  wire memDataQueue_io_deq_valid;
  wire[127:0] memDataQueue_io_deq_bits_data;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[135:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[4:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_2_io_out_bits_payload_manager_xact_id;
  wire LockingRRArbiter_2_io_out_bits_payload_uncached;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_g_type;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[25:0] LockingRRArbiter_3_io_out_bits_addr;
  wire[4:0] LockingRRArbiter_3_io_out_bits_tag;
  wire LockingRRArbiter_3_io_out_bits_rw;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[127:0] LockingRRArbiter_4_io_out_bits_data;
  wire LockingRRArbiter_5_io_in_0_ready;
  wire LockingRRArbiter_5_io_out_valid;
  wire LockingRRArbiter_5_io_out_bits_id;
  wire[16:0] LockingRRArbiter_5_io_out_bits_tag;
  wire[5:0] LockingRRArbiter_5_io_out_bits_idx;
  wire LockingRRArbiter_6_io_in_0_ready;
  wire LockingRRArbiter_6_io_out_valid;
  wire[16:0] LockingRRArbiter_6_io_out_bits_tag;
  wire[5:0] LockingRRArbiter_6_io_out_bits_idx;
  wire[7:0] LockingRRArbiter_6_io_out_bits_way_en;
  wire LockingRRArbiter_7_io_in_0_ready;
  wire LockingRRArbiter_7_io_out_valid;
  wire LockingRRArbiter_7_io_out_bits_id;
  wire[7:0] LockingRRArbiter_7_io_out_bits_addr;
  wire[7:0] LockingRRArbiter_7_io_out_bits_way_en;
  wire LockingRRArbiter_8_io_in_0_ready;
  wire LockingRRArbiter_8_io_out_valid;
  wire[127:0] LockingRRArbiter_8_io_out_bits_data;
  wire[7:0] LockingRRArbiter_8_io_out_bits_addr;
  wire[7:0] LockingRRArbiter_8_io_out_bits_way_en;
  wire[3:0] LockingRRArbiter_8_io_out_bits_wmask;


  assign T0 = acqQueue_io_deq_valid & T1;
  assign T1 = acq_conflict ^ 1'h1;
  assign acq_conflict = T2 != 1'h0;
  assign T2 = TagCacheTracker_io_acq_conflict;
  assign T3 = TagCacheTracker_io_uncached_acquire_ready & T4;
  assign T4 = acq_conflict ^ 1'h1;
  assign T5 = data_io_resp_valid & T6;
  assign T6 = 1'h0 == data_io_resp_bits_id;
  assign T7 = meta_io_resp_valid & T8;
  assign T8 = 1'h0 == meta_io_resp_bits_id;
  assign T9 = io_mem_resp_valid & T10;
  assign T10 = 4'h0 == T11;
  assign T11 = io_mem_resp_bits_tag >> 1'h1;
  assign T12 = acqQueue_io_deq_valid & T13;
  assign T13 = acq_conflict ^ 1'h1;
  assign io_mem_req_data_bits_data = memDataQueue_io_deq_bits_data;
  assign io_mem_req_data_valid = memDataQueue_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = memCMDQueue_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = memCMDQueue_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = memCMDQueue_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = memCMDQueue_io_deq_valid;
//  assign io_uncached_finish_ready = {1{$random}};
  assign io_uncached_grant_bits_payload_g_type = LockingRRArbiter_2_io_out_bits_payload_g_type;
  assign io_uncached_grant_bits_payload_uncached = LockingRRArbiter_2_io_out_bits_payload_uncached;
  assign io_uncached_grant_bits_payload_manager_xact_id = LockingRRArbiter_2_io_out_bits_payload_manager_xact_id;
  assign io_uncached_grant_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_uncached_grant_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_uncached_grant_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_uncached_grant_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_uncached_grant_valid = LockingRRArbiter_2_io_out_valid;
  assign io_uncached_acquire_ready = acqQueue_io_enq_ready;
  TagCacheMetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( LockingRRArbiter_5_io_out_valid ),
       .io_read_bits_id( LockingRRArbiter_5_io_out_bits_id ),
       .io_read_bits_tag( LockingRRArbiter_5_io_out_bits_tag ),
       .io_read_bits_idx( LockingRRArbiter_5_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( LockingRRArbiter_6_io_out_valid ),
       .io_write_bits_tag( LockingRRArbiter_6_io_out_bits_tag ),
       .io_write_bits_idx( LockingRRArbiter_6_io_out_bits_idx ),
       .io_write_bits_way_en( LockingRRArbiter_6_io_out_bits_way_en ),
       .io_resp_valid( meta_io_resp_valid ),
       .io_resp_bits_id( meta_io_resp_bits_id ),
       .io_resp_bits_tag( meta_io_resp_bits_tag ),
       .io_resp_bits_hit( meta_io_resp_bits_hit ),
       .io_resp_bits_way_en( meta_io_resp_bits_way_en )
  );
  TagCacheDataArray data(.clk(clk),
       .io_read_ready( data_io_read_ready ),
       .io_read_valid( LockingRRArbiter_7_io_out_valid ),
       .io_read_bits_id( LockingRRArbiter_7_io_out_bits_id ),
       .io_read_bits_addr( LockingRRArbiter_7_io_out_bits_addr ),
       .io_read_bits_way_en( LockingRRArbiter_7_io_out_bits_way_en ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( LockingRRArbiter_8_io_out_valid ),
       .io_write_bits_data( LockingRRArbiter_8_io_out_bits_data ),
       .io_write_bits_addr( LockingRRArbiter_8_io_out_bits_addr ),
       .io_write_bits_way_en( LockingRRArbiter_8_io_out_bits_way_en ),
       .io_write_bits_wmask( LockingRRArbiter_8_io_out_bits_wmask ),
       .io_resp_valid( data_io_resp_valid ),
       .io_resp_bits_id( data_io_resp_bits_id ),
       .io_resp_bits_data( data_io_resp_bits_data )
  );
  TagCacheTracker TagCacheTracker(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( TagCacheTracker_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( T12 ),
       .io_uncached_acquire_bits_header_src( acqQueue_io_deq_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( acqQueue_io_deq_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( acqQueue_io_deq_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( acqQueue_io_deq_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( acqQueue_io_deq_bits_payload_data ),
       .io_uncached_acquire_bits_payload_uncached( acqQueue_io_deq_bits_payload_uncached ),
       .io_uncached_acquire_bits_payload_a_type( acqQueue_io_deq_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_subblock( acqQueue_io_deq_bits_payload_subblock ),
       .io_uncached_grant_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_uncached_grant_valid( TagCacheTracker_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( TagCacheTracker_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( TagCacheTracker_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_manager_xact_id( TagCacheTracker_io_uncached_grant_bits_payload_manager_xact_id ),
       .io_uncached_grant_bits_payload_uncached( TagCacheTracker_io_uncached_grant_bits_payload_uncached ),
       .io_uncached_grant_bits_payload_g_type( TagCacheTracker_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       //.io_uncached_finish_valid(  )
       //.io_uncached_finish_bits_header_src(  )
       //.io_uncached_finish_bits_header_dst(  )
       //.io_uncached_finish_bits_payload_manager_xact_id(  )
       .io_mem_req_cmd_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_mem_req_cmd_valid( TagCacheTracker_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( TagCacheTracker_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( TagCacheTracker_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( TagCacheTracker_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_mem_req_data_valid( TagCacheTracker_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( TagCacheTracker_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( T9 ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_meta_read_ready( LockingRRArbiter_5_io_in_0_ready ),
       .io_meta_read_valid( TagCacheTracker_io_meta_read_valid ),
       .io_meta_read_bits_id( TagCacheTracker_io_meta_read_bits_id ),
       .io_meta_read_bits_tag( TagCacheTracker_io_meta_read_bits_tag ),
       .io_meta_read_bits_idx( TagCacheTracker_io_meta_read_bits_idx ),
       .io_meta_write_ready( LockingRRArbiter_6_io_in_0_ready ),
       .io_meta_write_valid( TagCacheTracker_io_meta_write_valid ),
       .io_meta_write_bits_tag( TagCacheTracker_io_meta_write_bits_tag ),
       .io_meta_write_bits_idx( TagCacheTracker_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( TagCacheTracker_io_meta_write_bits_way_en ),
       .io_meta_resp_valid( T7 ),
       .io_meta_resp_bits_id( meta_io_resp_bits_id ),
       .io_meta_resp_bits_tag( meta_io_resp_bits_tag ),
       .io_meta_resp_bits_hit( meta_io_resp_bits_hit ),
       .io_meta_resp_bits_way_en( meta_io_resp_bits_way_en ),
       .io_data_read_ready( LockingRRArbiter_7_io_in_0_ready ),
       .io_data_read_valid( TagCacheTracker_io_data_read_valid ),
       .io_data_read_bits_id( TagCacheTracker_io_data_read_bits_id ),
       .io_data_read_bits_addr( TagCacheTracker_io_data_read_bits_addr ),
       .io_data_read_bits_way_en( TagCacheTracker_io_data_read_bits_way_en ),
       .io_data_write_ready( LockingRRArbiter_8_io_in_0_ready ),
       .io_data_write_valid( TagCacheTracker_io_data_write_valid ),
       .io_data_write_bits_data( TagCacheTracker_io_data_write_bits_data ),
       .io_data_write_bits_addr( TagCacheTracker_io_data_write_bits_addr ),
       .io_data_write_bits_way_en( TagCacheTracker_io_data_write_bits_way_en ),
       .io_data_write_bits_wmask( TagCacheTracker_io_data_write_bits_wmask ),
       .io_data_resp_valid( T5 ),
       .io_data_resp_bits_id( data_io_resp_bits_id ),
       .io_data_resp_bits_data( data_io_resp_bits_data ),
       .io_acq_conflict( TagCacheTracker_io_acq_conflict )
       //.io_acq_match(  )
  );
  Queue_9 acqQueue(.clk(clk), .reset(reset),
       .io_enq_ready( acqQueue_io_enq_ready ),
       .io_enq_valid( io_uncached_acquire_valid ),
       .io_enq_bits_header_src( io_uncached_acquire_bits_header_src ),
       .io_enq_bits_header_dst( io_uncached_acquire_bits_header_dst ),
       .io_enq_bits_payload_addr( io_uncached_acquire_bits_payload_addr ),
       .io_enq_bits_payload_client_xact_id( io_uncached_acquire_bits_payload_client_xact_id ),
       .io_enq_bits_payload_data( io_uncached_acquire_bits_payload_data ),
       .io_enq_bits_payload_uncached( io_uncached_acquire_bits_payload_uncached ),
       .io_enq_bits_payload_a_type( io_uncached_acquire_bits_payload_a_type ),
       .io_enq_bits_payload_subblock( io_uncached_acquire_bits_payload_subblock ),
       .io_deq_ready( T3 ),
       .io_deq_valid( acqQueue_io_deq_valid ),
       .io_deq_bits_header_src( acqQueue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( acqQueue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( acqQueue_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( acqQueue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( acqQueue_io_deq_bits_payload_data ),
       .io_deq_bits_payload_uncached( acqQueue_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_a_type( acqQueue_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_subblock( acqQueue_io_deq_bits_payload_subblock )
       //.io_count(  )
  );
  Queue_10 memCMDQueue(.clk(clk), .reset(reset),
       .io_enq_ready( memCMDQueue_io_enq_ready ),
       .io_enq_valid( LockingRRArbiter_3_io_out_valid ),
       .io_enq_bits_addr( LockingRRArbiter_3_io_out_bits_addr ),
       .io_enq_bits_tag( LockingRRArbiter_3_io_out_bits_tag ),
       .io_enq_bits_rw( LockingRRArbiter_3_io_out_bits_rw ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( memCMDQueue_io_deq_valid ),
       .io_deq_bits_addr( memCMDQueue_io_deq_bits_addr ),
       .io_deq_bits_tag( memCMDQueue_io_deq_bits_tag ),
       .io_deq_bits_rw( memCMDQueue_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_11 memDataQueue(.clk(clk), .reset(reset),
       .io_enq_ready( memDataQueue_io_enq_ready ),
       .io_enq_valid( LockingRRArbiter_4_io_out_valid ),
       .io_enq_bits_data( LockingRRArbiter_4_io_out_bits_data ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( memDataQueue_io_deq_valid ),
       .io_deq_bits_data( memDataQueue_io_deq_bits_data )
       //.io_count(  )
  );
  Arbiter_11 acq_arb(
       //.io_in_0_ready(  )
       .io_in_0_valid( TagCacheTracker_io_uncached_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T0 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign acq_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  LockingRRArbiter_2 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_uncached_grant_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       .io_in_0_bits_payload_data( TagCacheTracker_io_uncached_grant_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( TagCacheTracker_io_uncached_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_manager_xact_id( TagCacheTracker_io_uncached_grant_bits_payload_manager_xact_id ),
       .io_in_0_bits_payload_uncached( TagCacheTracker_io_uncached_grant_bits_payload_uncached ),
       .io_in_0_bits_payload_g_type( TagCacheTracker_io_uncached_grant_bits_payload_g_type ),
       .io_out_ready( io_uncached_grant_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_manager_xact_id( LockingRRArbiter_2_io_out_bits_payload_manager_xact_id ),
       .io_out_bits_payload_uncached( LockingRRArbiter_2_io_out_bits_payload_uncached ),
       .io_out_bits_payload_g_type( LockingRRArbiter_2_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign LockingRRArbiter_2.io_in_0_bits_header_src = {1{$random}};
    assign LockingRRArbiter_2.io_in_0_bits_header_dst = {1{$random}};
// synthesis translate_on
`endif
  LockingRRArbiter_3 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_mem_req_cmd_valid ),
       .io_in_0_bits_addr( TagCacheTracker_io_mem_req_cmd_bits_addr ),
       .io_in_0_bits_tag( TagCacheTracker_io_mem_req_cmd_bits_tag ),
       .io_in_0_bits_rw( TagCacheTracker_io_mem_req_cmd_bits_rw ),
       .io_out_ready( memCMDQueue_io_enq_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_addr( LockingRRArbiter_3_io_out_bits_addr ),
       .io_out_bits_tag( LockingRRArbiter_3_io_out_bits_tag ),
       .io_out_bits_rw( LockingRRArbiter_3_io_out_bits_rw )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_mem_req_data_valid ),
       .io_in_0_bits_data( TagCacheTracker_io_mem_req_data_bits_data ),
       .io_out_ready( memDataQueue_io_enq_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_data( LockingRRArbiter_4_io_out_bits_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_5 LockingRRArbiter_5(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_5_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_meta_read_valid ),
       .io_in_0_bits_id( TagCacheTracker_io_meta_read_bits_id ),
       .io_in_0_bits_tag( TagCacheTracker_io_meta_read_bits_tag ),
       .io_in_0_bits_idx( TagCacheTracker_io_meta_read_bits_idx ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( LockingRRArbiter_5_io_out_valid ),
       .io_out_bits_id( LockingRRArbiter_5_io_out_bits_id ),
       .io_out_bits_tag( LockingRRArbiter_5_io_out_bits_tag ),
       .io_out_bits_idx( LockingRRArbiter_5_io_out_bits_idx )
       //.io_chosen(  )
  );
  LockingRRArbiter_6 LockingRRArbiter_6(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_6_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_meta_write_valid ),
       .io_in_0_bits_tag( TagCacheTracker_io_meta_write_bits_tag ),
       .io_in_0_bits_idx( TagCacheTracker_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( TagCacheTracker_io_meta_write_bits_way_en ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( LockingRRArbiter_6_io_out_valid ),
       .io_out_bits_tag( LockingRRArbiter_6_io_out_bits_tag ),
       .io_out_bits_idx( LockingRRArbiter_6_io_out_bits_idx ),
       .io_out_bits_way_en( LockingRRArbiter_6_io_out_bits_way_en )
       //.io_chosen(  )
  );
  LockingRRArbiter_7 LockingRRArbiter_7(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_7_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_data_read_valid ),
       .io_in_0_bits_id( TagCacheTracker_io_data_read_bits_id ),
       .io_in_0_bits_addr( TagCacheTracker_io_data_read_bits_addr ),
       .io_in_0_bits_way_en( TagCacheTracker_io_data_read_bits_way_en ),
       .io_out_ready( data_io_read_ready ),
       .io_out_valid( LockingRRArbiter_7_io_out_valid ),
       .io_out_bits_id( LockingRRArbiter_7_io_out_bits_id ),
       .io_out_bits_addr( LockingRRArbiter_7_io_out_bits_addr ),
       .io_out_bits_way_en( LockingRRArbiter_7_io_out_bits_way_en )
       //.io_chosen(  )
  );
  LockingRRArbiter_8 LockingRRArbiter_8(.clk(clk), .reset(reset),
       .io_in_0_ready( LockingRRArbiter_8_io_in_0_ready ),
       .io_in_0_valid( TagCacheTracker_io_data_write_valid ),
       .io_in_0_bits_data( TagCacheTracker_io_data_write_bits_data ),
       .io_in_0_bits_addr( TagCacheTracker_io_data_write_bits_addr ),
       .io_in_0_bits_way_en( TagCacheTracker_io_data_write_bits_way_en ),
       .io_in_0_bits_wmask( TagCacheTracker_io_data_write_bits_wmask ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( LockingRRArbiter_8_io_out_valid ),
       .io_out_bits_data( LockingRRArbiter_8_io_out_bits_data ),
       .io_out_bits_addr( LockingRRArbiter_8_io_out_bits_addr ),
       .io_out_bits_way_en( LockingRRArbiter_8_io_out_bits_way_en ),
       .io_out_bits_wmask( LockingRRArbiter_8_io_out_bits_wmask )
       //.io_chosen(  )
  );
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [135:0] io_tiles_0_acquire_bits_payload_data,
    input  io_tiles_0_acquire_bits_payload_uncached,
    input [1:0] io_tiles_0_acquire_bits_payload_a_type,
    input [128:0] io_tiles_0_acquire_bits_payload_subblock,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[135:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_manager_xact_id,
    output io_tiles_0_grant_bits_payload_uncached,
    output[1:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [3:0] io_tiles_0_finish_bits_payload_manager_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [135:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_acquire_ready,
    input  io_htif_acquire_valid,
    input [1:0] io_htif_acquire_bits_header_src,
    input [1:0] io_htif_acquire_bits_header_dst,
    input [25:0] io_htif_acquire_bits_payload_addr,
    input [1:0] io_htif_acquire_bits_payload_client_xact_id,
    input [135:0] io_htif_acquire_bits_payload_data,
    input  io_htif_acquire_bits_payload_uncached,
    input [1:0] io_htif_acquire_bits_payload_a_type,
    input [128:0] io_htif_acquire_bits_payload_subblock,
    input  io_htif_grant_ready,
    output io_htif_grant_valid,
    output[1:0] io_htif_grant_bits_header_src,
    output[1:0] io_htif_grant_bits_header_dst,
    output[135:0] io_htif_grant_bits_payload_data,
    output[1:0] io_htif_grant_bits_payload_client_xact_id,
    output[3:0] io_htif_grant_bits_payload_manager_xact_id,
    output io_htif_grant_bits_payload_uncached,
    output[1:0] io_htif_grant_bits_payload_g_type,
    output io_htif_finish_ready,
    input  io_htif_finish_valid,
    input [1:0] io_htif_finish_bits_header_src,
    input [1:0] io_htif_finish_bits_header_dst,
    input [3:0] io_htif_finish_bits_payload_manager_xact_id,
    input  io_htif_probe_ready,
    output io_htif_probe_valid,
    output[1:0] io_htif_probe_bits_header_src,
    output[1:0] io_htif_probe_bits_header_dst,
    output[25:0] io_htif_probe_bits_payload_addr,
    output[1:0] io_htif_probe_bits_payload_p_type,
    output io_htif_release_ready,
    input  io_htif_release_valid,
    input [1:0] io_htif_release_bits_header_src,
    input [1:0] io_htif_release_bits_header_dst,
    input [25:0] io_htif_release_bits_payload_addr,
    input [1:0] io_htif_release_bits_payload_client_xact_id,
    input [135:0] io_htif_release_bits_payload_data,
    input [2:0] io_htif_release_bits_payload_r_type,
    input  io_incoherent_1,
    input  io_incoherent_0,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire tagCache_io_uncached_acquire_ready;
  wire tagCache_io_uncached_grant_valid;
  wire[1:0] tagCache_io_uncached_grant_bits_header_src;
  wire[1:0] tagCache_io_uncached_grant_bits_header_dst;
  wire[135:0] tagCache_io_uncached_grant_bits_payload_data;
  wire[4:0] tagCache_io_uncached_grant_bits_payload_client_xact_id;
  wire tagCache_io_uncached_grant_bits_payload_manager_xact_id;
  wire tagCache_io_uncached_grant_bits_payload_uncached;
  wire[1:0] tagCache_io_uncached_grant_bits_payload_g_type;
  wire tagCache_io_mem_req_cmd_valid;
  wire[25:0] tagCache_io_mem_req_cmd_bits_addr;
  wire[4:0] tagCache_io_mem_req_cmd_bits_tag;
  wire tagCache_io_mem_req_cmd_bits_rw;
  wire tagCache_io_mem_req_data_valid;
  wire[127:0] tagCache_io_mem_req_data_bits_data;
  wire net_io_clients_1_acquire_ready;
  wire net_io_clients_1_grant_valid;
  wire[1:0] net_io_clients_1_grant_bits_header_src;
  wire[1:0] net_io_clients_1_grant_bits_header_dst;
  wire[135:0] net_io_clients_1_grant_bits_payload_data;
  wire[1:0] net_io_clients_1_grant_bits_payload_client_xact_id;
  wire[3:0] net_io_clients_1_grant_bits_payload_manager_xact_id;
  wire net_io_clients_1_grant_bits_payload_uncached;
  wire[1:0] net_io_clients_1_grant_bits_payload_g_type;
  wire net_io_clients_1_finish_ready;
  wire net_io_clients_1_probe_valid;
  wire[1:0] net_io_clients_1_probe_bits_header_src;
  wire[1:0] net_io_clients_1_probe_bits_header_dst;
  wire[25:0] net_io_clients_1_probe_bits_payload_addr;
  wire[1:0] net_io_clients_1_probe_bits_payload_p_type;
  wire net_io_clients_1_release_ready;
  wire net_io_clients_0_acquire_ready;
  wire net_io_clients_0_grant_valid;
  wire[1:0] net_io_clients_0_grant_bits_header_src;
  wire[1:0] net_io_clients_0_grant_bits_header_dst;
  wire[135:0] net_io_clients_0_grant_bits_payload_data;
  wire[1:0] net_io_clients_0_grant_bits_payload_client_xact_id;
  wire[3:0] net_io_clients_0_grant_bits_payload_manager_xact_id;
  wire net_io_clients_0_grant_bits_payload_uncached;
  wire[1:0] net_io_clients_0_grant_bits_payload_g_type;
  wire net_io_clients_0_finish_ready;
  wire net_io_clients_0_probe_valid;
  wire[1:0] net_io_clients_0_probe_bits_header_src;
  wire[1:0] net_io_clients_0_probe_bits_header_dst;
  wire[25:0] net_io_clients_0_probe_bits_payload_addr;
  wire[1:0] net_io_clients_0_probe_bits_payload_p_type;
  wire net_io_clients_0_release_ready;
  wire net_io_managers_0_acquire_valid;
  wire[1:0] net_io_managers_0_acquire_bits_header_src;
  wire[1:0] net_io_managers_0_acquire_bits_header_dst;
  wire[25:0] net_io_managers_0_acquire_bits_payload_addr;
  wire[1:0] net_io_managers_0_acquire_bits_payload_client_xact_id;
  wire[135:0] net_io_managers_0_acquire_bits_payload_data;
  wire net_io_managers_0_acquire_bits_payload_uncached;
  wire[1:0] net_io_managers_0_acquire_bits_payload_a_type;
  wire[128:0] net_io_managers_0_acquire_bits_payload_subblock;
  wire net_io_managers_0_grant_ready;
  wire net_io_managers_0_finish_valid;
  wire[1:0] net_io_managers_0_finish_bits_header_src;
  wire[1:0] net_io_managers_0_finish_bits_header_dst;
  wire[3:0] net_io_managers_0_finish_bits_payload_manager_xact_id;
  wire net_io_managers_0_probe_ready;
  wire net_io_managers_0_release_valid;
  wire[1:0] net_io_managers_0_release_bits_header_src;
  wire[1:0] net_io_managers_0_release_bits_header_dst;
  wire[25:0] net_io_managers_0_release_bits_payload_addr;
  wire[1:0] net_io_managers_0_release_bits_payload_client_xact_id;
  wire[135:0] net_io_managers_0_release_bits_payload_data;
  wire[2:0] net_io_managers_0_release_bits_payload_r_type;
  wire L2BroadcastHub_io_inner_acquire_ready;
  wire L2BroadcastHub_io_inner_grant_valid;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_header_src;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_header_dst;
  wire[135:0] L2BroadcastHub_io_inner_grant_bits_payload_data;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_payload_client_xact_id;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_payload_manager_xact_id;
  wire L2BroadcastHub_io_inner_grant_bits_payload_uncached;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_payload_g_type;
  wire L2BroadcastHub_io_inner_finish_ready;
  wire L2BroadcastHub_io_inner_probe_valid;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_header_src;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_header_dst;
  wire[25:0] L2BroadcastHub_io_inner_probe_bits_payload_addr;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_payload_p_type;
  wire L2BroadcastHub_io_inner_release_ready;
  wire L2BroadcastHub_io_outer_acquire_valid;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_header_src;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_header_dst;
  wire[25:0] L2BroadcastHub_io_outer_acquire_bits_payload_addr;
  wire[4:0] L2BroadcastHub_io_outer_acquire_bits_payload_client_xact_id;
  wire[135:0] L2BroadcastHub_io_outer_acquire_bits_payload_data;
  wire L2BroadcastHub_io_outer_acquire_bits_payload_uncached;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_payload_a_type;
  wire[128:0] L2BroadcastHub_io_outer_acquire_bits_payload_subblock;
  wire L2BroadcastHub_io_outer_grant_ready;
  wire L2BroadcastHub_io_outer_finish_valid;
  wire[1:0] L2BroadcastHub_io_outer_finish_bits_header_src;
  wire[1:0] L2BroadcastHub_io_outer_finish_bits_header_dst;
  wire L2BroadcastHub_io_outer_finish_bits_payload_manager_xact_id;


//  assign io_mem_backup_req_bits = {1{$random}};
//  assign io_mem_backup_req_valid = {1{$random}};
//  assign io_mem_resp_ready = {1{$random}};
  assign io_mem_req_data_bits_data = tagCache_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = tagCache_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = tagCache_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = tagCache_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = tagCache_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = tagCache_io_mem_req_cmd_valid;
  assign io_htif_release_ready = net_io_clients_1_release_ready;
  assign io_htif_probe_bits_payload_p_type = net_io_clients_1_probe_bits_payload_p_type;
  assign io_htif_probe_bits_payload_addr = net_io_clients_1_probe_bits_payload_addr;
  assign io_htif_probe_bits_header_dst = net_io_clients_1_probe_bits_header_dst;
  assign io_htif_probe_bits_header_src = net_io_clients_1_probe_bits_header_src;
  assign io_htif_probe_valid = net_io_clients_1_probe_valid;
  assign io_htif_finish_ready = net_io_clients_1_finish_ready;
  assign io_htif_grant_bits_payload_g_type = net_io_clients_1_grant_bits_payload_g_type;
  assign io_htif_grant_bits_payload_uncached = net_io_clients_1_grant_bits_payload_uncached;
  assign io_htif_grant_bits_payload_manager_xact_id = net_io_clients_1_grant_bits_payload_manager_xact_id;
  assign io_htif_grant_bits_payload_client_xact_id = net_io_clients_1_grant_bits_payload_client_xact_id;
  assign io_htif_grant_bits_payload_data = net_io_clients_1_grant_bits_payload_data;
  assign io_htif_grant_bits_header_dst = net_io_clients_1_grant_bits_header_dst;
  assign io_htif_grant_bits_header_src = net_io_clients_1_grant_bits_header_src;
  assign io_htif_grant_valid = net_io_clients_1_grant_valid;
  assign io_htif_acquire_ready = net_io_clients_1_acquire_ready;
  assign io_tiles_0_release_ready = net_io_clients_0_release_ready;
  assign io_tiles_0_probe_bits_payload_p_type = net_io_clients_0_probe_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_addr = net_io_clients_0_probe_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = net_io_clients_0_probe_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = net_io_clients_0_probe_bits_header_src;
  assign io_tiles_0_probe_valid = net_io_clients_0_probe_valid;
  assign io_tiles_0_finish_ready = net_io_clients_0_finish_ready;
  assign io_tiles_0_grant_bits_payload_g_type = net_io_clients_0_grant_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_uncached = net_io_clients_0_grant_bits_payload_uncached;
  assign io_tiles_0_grant_bits_payload_manager_xact_id = net_io_clients_0_grant_bits_payload_manager_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = net_io_clients_0_grant_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = net_io_clients_0_grant_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = net_io_clients_0_grant_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = net_io_clients_0_grant_bits_header_src;
  assign io_tiles_0_grant_valid = net_io_clients_0_grant_valid;
  assign io_tiles_0_acquire_ready = net_io_clients_0_acquire_ready;
  RocketChipCrossbarNetwork net(.clk(clk), .reset(reset),
       .io_clients_1_acquire_ready( net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( io_htif_acquire_valid ),
       .io_clients_1_acquire_bits_header_src( io_htif_acquire_bits_header_src ),
       .io_clients_1_acquire_bits_header_dst( io_htif_acquire_bits_header_dst ),
       .io_clients_1_acquire_bits_payload_addr( io_htif_acquire_bits_payload_addr ),
       .io_clients_1_acquire_bits_payload_client_xact_id( io_htif_acquire_bits_payload_client_xact_id ),
       .io_clients_1_acquire_bits_payload_data( io_htif_acquire_bits_payload_data ),
       .io_clients_1_acquire_bits_payload_uncached( io_htif_acquire_bits_payload_uncached ),
       .io_clients_1_acquire_bits_payload_a_type( io_htif_acquire_bits_payload_a_type ),
       .io_clients_1_acquire_bits_payload_subblock( io_htif_acquire_bits_payload_subblock ),
       .io_clients_1_grant_ready( io_htif_grant_ready ),
       .io_clients_1_grant_valid( net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_header_src( net_io_clients_1_grant_bits_header_src ),
       .io_clients_1_grant_bits_header_dst( net_io_clients_1_grant_bits_header_dst ),
       .io_clients_1_grant_bits_payload_data( net_io_clients_1_grant_bits_payload_data ),
       .io_clients_1_grant_bits_payload_client_xact_id( net_io_clients_1_grant_bits_payload_client_xact_id ),
       .io_clients_1_grant_bits_payload_manager_xact_id( net_io_clients_1_grant_bits_payload_manager_xact_id ),
       .io_clients_1_grant_bits_payload_uncached( net_io_clients_1_grant_bits_payload_uncached ),
       .io_clients_1_grant_bits_payload_g_type( net_io_clients_1_grant_bits_payload_g_type ),
       .io_clients_1_finish_ready( net_io_clients_1_finish_ready ),
       .io_clients_1_finish_valid( io_htif_finish_valid ),
       .io_clients_1_finish_bits_header_src( io_htif_finish_bits_header_src ),
       .io_clients_1_finish_bits_header_dst( io_htif_finish_bits_header_dst ),
       .io_clients_1_finish_bits_payload_manager_xact_id( io_htif_finish_bits_payload_manager_xact_id ),
       .io_clients_1_probe_ready( io_htif_probe_ready ),
       .io_clients_1_probe_valid( net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_header_src( net_io_clients_1_probe_bits_header_src ),
       .io_clients_1_probe_bits_header_dst( net_io_clients_1_probe_bits_header_dst ),
       .io_clients_1_probe_bits_payload_addr( net_io_clients_1_probe_bits_payload_addr ),
       .io_clients_1_probe_bits_payload_p_type( net_io_clients_1_probe_bits_payload_p_type ),
       .io_clients_1_release_ready( net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( io_htif_release_valid ),
       .io_clients_1_release_bits_header_src( io_htif_release_bits_header_src ),
       .io_clients_1_release_bits_header_dst( io_htif_release_bits_header_dst ),
       .io_clients_1_release_bits_payload_addr( io_htif_release_bits_payload_addr ),
       .io_clients_1_release_bits_payload_client_xact_id( io_htif_release_bits_payload_client_xact_id ),
       .io_clients_1_release_bits_payload_data( io_htif_release_bits_payload_data ),
       .io_clients_1_release_bits_payload_r_type( io_htif_release_bits_payload_r_type ),
       .io_clients_0_acquire_ready( net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_0_acquire_valid ),
       .io_clients_0_acquire_bits_header_src( io_tiles_0_acquire_bits_header_src ),
       .io_clients_0_acquire_bits_header_dst( io_tiles_0_acquire_bits_header_dst ),
       .io_clients_0_acquire_bits_payload_addr( io_tiles_0_acquire_bits_payload_addr ),
       .io_clients_0_acquire_bits_payload_client_xact_id( io_tiles_0_acquire_bits_payload_client_xact_id ),
       .io_clients_0_acquire_bits_payload_data( io_tiles_0_acquire_bits_payload_data ),
       .io_clients_0_acquire_bits_payload_uncached( io_tiles_0_acquire_bits_payload_uncached ),
       .io_clients_0_acquire_bits_payload_a_type( io_tiles_0_acquire_bits_payload_a_type ),
       .io_clients_0_acquire_bits_payload_subblock( io_tiles_0_acquire_bits_payload_subblock ),
       .io_clients_0_grant_ready( io_tiles_0_grant_ready ),
       .io_clients_0_grant_valid( net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_header_src( net_io_clients_0_grant_bits_header_src ),
       .io_clients_0_grant_bits_header_dst( net_io_clients_0_grant_bits_header_dst ),
       .io_clients_0_grant_bits_payload_data( net_io_clients_0_grant_bits_payload_data ),
       .io_clients_0_grant_bits_payload_client_xact_id( net_io_clients_0_grant_bits_payload_client_xact_id ),
       .io_clients_0_grant_bits_payload_manager_xact_id( net_io_clients_0_grant_bits_payload_manager_xact_id ),
       .io_clients_0_grant_bits_payload_uncached( net_io_clients_0_grant_bits_payload_uncached ),
       .io_clients_0_grant_bits_payload_g_type( net_io_clients_0_grant_bits_payload_g_type ),
       .io_clients_0_finish_ready( net_io_clients_0_finish_ready ),
       .io_clients_0_finish_valid( io_tiles_0_finish_valid ),
       .io_clients_0_finish_bits_header_src( io_tiles_0_finish_bits_header_src ),
       .io_clients_0_finish_bits_header_dst( io_tiles_0_finish_bits_header_dst ),
       .io_clients_0_finish_bits_payload_manager_xact_id( io_tiles_0_finish_bits_payload_manager_xact_id ),
       .io_clients_0_probe_ready( io_tiles_0_probe_ready ),
       .io_clients_0_probe_valid( net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_header_src( net_io_clients_0_probe_bits_header_src ),
       .io_clients_0_probe_bits_header_dst( net_io_clients_0_probe_bits_header_dst ),
       .io_clients_0_probe_bits_payload_addr( net_io_clients_0_probe_bits_payload_addr ),
       .io_clients_0_probe_bits_payload_p_type( net_io_clients_0_probe_bits_payload_p_type ),
       .io_clients_0_release_ready( net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_0_release_valid ),
       .io_clients_0_release_bits_header_src( io_tiles_0_release_bits_header_src ),
       .io_clients_0_release_bits_header_dst( io_tiles_0_release_bits_header_dst ),
       .io_clients_0_release_bits_payload_addr( io_tiles_0_release_bits_payload_addr ),
       .io_clients_0_release_bits_payload_client_xact_id( io_tiles_0_release_bits_payload_client_xact_id ),
       .io_clients_0_release_bits_payload_data( io_tiles_0_release_bits_payload_data ),
       .io_clients_0_release_bits_payload_r_type( io_tiles_0_release_bits_payload_r_type ),
       .io_managers_0_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_managers_0_acquire_valid( net_io_managers_0_acquire_valid ),
       .io_managers_0_acquire_bits_header_src( net_io_managers_0_acquire_bits_header_src ),
       .io_managers_0_acquire_bits_header_dst( net_io_managers_0_acquire_bits_header_dst ),
       .io_managers_0_acquire_bits_payload_addr( net_io_managers_0_acquire_bits_payload_addr ),
       .io_managers_0_acquire_bits_payload_client_xact_id( net_io_managers_0_acquire_bits_payload_client_xact_id ),
       .io_managers_0_acquire_bits_payload_data( net_io_managers_0_acquire_bits_payload_data ),
       .io_managers_0_acquire_bits_payload_uncached( net_io_managers_0_acquire_bits_payload_uncached ),
       .io_managers_0_acquire_bits_payload_a_type( net_io_managers_0_acquire_bits_payload_a_type ),
       .io_managers_0_acquire_bits_payload_subblock( net_io_managers_0_acquire_bits_payload_subblock ),
       .io_managers_0_grant_ready( net_io_managers_0_grant_ready ),
       .io_managers_0_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_managers_0_grant_bits_header_src( L2BroadcastHub_io_inner_grant_bits_header_src ),
       .io_managers_0_grant_bits_header_dst( L2BroadcastHub_io_inner_grant_bits_header_dst ),
       .io_managers_0_grant_bits_payload_data( L2BroadcastHub_io_inner_grant_bits_payload_data ),
       .io_managers_0_grant_bits_payload_client_xact_id( L2BroadcastHub_io_inner_grant_bits_payload_client_xact_id ),
       .io_managers_0_grant_bits_payload_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_payload_manager_xact_id ),
       .io_managers_0_grant_bits_payload_uncached( L2BroadcastHub_io_inner_grant_bits_payload_uncached ),
       .io_managers_0_grant_bits_payload_g_type( L2BroadcastHub_io_inner_grant_bits_payload_g_type ),
       .io_managers_0_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_managers_0_finish_valid( net_io_managers_0_finish_valid ),
       .io_managers_0_finish_bits_header_src( net_io_managers_0_finish_bits_header_src ),
       .io_managers_0_finish_bits_header_dst( net_io_managers_0_finish_bits_header_dst ),
       .io_managers_0_finish_bits_payload_manager_xact_id( net_io_managers_0_finish_bits_payload_manager_xact_id ),
       .io_managers_0_probe_ready( net_io_managers_0_probe_ready ),
       .io_managers_0_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_managers_0_probe_bits_header_src( L2BroadcastHub_io_inner_probe_bits_header_src ),
       .io_managers_0_probe_bits_header_dst( L2BroadcastHub_io_inner_probe_bits_header_dst ),
       .io_managers_0_probe_bits_payload_addr( L2BroadcastHub_io_inner_probe_bits_payload_addr ),
       .io_managers_0_probe_bits_payload_p_type( L2BroadcastHub_io_inner_probe_bits_payload_p_type ),
       .io_managers_0_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_managers_0_release_valid( net_io_managers_0_release_valid ),
       .io_managers_0_release_bits_header_src( net_io_managers_0_release_bits_header_src ),
       .io_managers_0_release_bits_header_dst( net_io_managers_0_release_bits_header_dst ),
       .io_managers_0_release_bits_payload_addr( net_io_managers_0_release_bits_payload_addr ),
       .io_managers_0_release_bits_payload_client_xact_id( net_io_managers_0_release_bits_payload_client_xact_id ),
       .io_managers_0_release_bits_payload_data( net_io_managers_0_release_bits_payload_data ),
       .io_managers_0_release_bits_payload_r_type( net_io_managers_0_release_bits_payload_r_type )
  );
  L2BroadcastHub L2BroadcastHub(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_inner_acquire_valid( net_io_managers_0_acquire_valid ),
       .io_inner_acquire_bits_header_src( net_io_managers_0_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( net_io_managers_0_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( net_io_managers_0_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( net_io_managers_0_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( net_io_managers_0_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_uncached( net_io_managers_0_acquire_bits_payload_uncached ),
       .io_inner_acquire_bits_payload_a_type( net_io_managers_0_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_subblock( net_io_managers_0_acquire_bits_payload_subblock ),
       .io_inner_grant_ready( net_io_managers_0_grant_ready ),
       .io_inner_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( L2BroadcastHub_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( L2BroadcastHub_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( L2BroadcastHub_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( L2BroadcastHub_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_payload_manager_xact_id ),
       .io_inner_grant_bits_payload_uncached( L2BroadcastHub_io_inner_grant_bits_payload_uncached ),
       .io_inner_grant_bits_payload_g_type( L2BroadcastHub_io_inner_grant_bits_payload_g_type ),
       .io_inner_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_inner_finish_valid( net_io_managers_0_finish_valid ),
       .io_inner_finish_bits_header_src( net_io_managers_0_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( net_io_managers_0_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_manager_xact_id( net_io_managers_0_finish_bits_payload_manager_xact_id ),
       .io_inner_probe_ready( net_io_managers_0_probe_ready ),
       .io_inner_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( L2BroadcastHub_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( L2BroadcastHub_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( L2BroadcastHub_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_p_type( L2BroadcastHub_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_inner_release_valid( net_io_managers_0_release_valid ),
       .io_inner_release_bits_header_src( net_io_managers_0_release_bits_header_src ),
       .io_inner_release_bits_header_dst( net_io_managers_0_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( net_io_managers_0_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( net_io_managers_0_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_data( net_io_managers_0_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( net_io_managers_0_release_bits_payload_r_type ),
       .io_outer_acquire_ready( tagCache_io_uncached_acquire_ready ),
       .io_outer_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( L2BroadcastHub_io_outer_acquire_bits_header_src ),
       .io_outer_acquire_bits_header_dst( L2BroadcastHub_io_outer_acquire_bits_header_dst ),
       .io_outer_acquire_bits_payload_addr( L2BroadcastHub_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( L2BroadcastHub_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_uncached( L2BroadcastHub_io_outer_acquire_bits_payload_uncached ),
       .io_outer_acquire_bits_payload_a_type( L2BroadcastHub_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_subblock( L2BroadcastHub_io_outer_acquire_bits_payload_subblock ),
       .io_outer_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_outer_grant_valid( tagCache_io_uncached_grant_valid ),
       .io_outer_grant_bits_header_src( tagCache_io_uncached_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( tagCache_io_uncached_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( tagCache_io_uncached_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( tagCache_io_uncached_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_manager_xact_id( tagCache_io_uncached_grant_bits_payload_manager_xact_id ),
       .io_outer_grant_bits_payload_uncached( tagCache_io_uncached_grant_bits_payload_uncached ),
       .io_outer_grant_bits_payload_g_type( tagCache_io_uncached_grant_bits_payload_g_type ),
       //.io_outer_finish_ready(  )
       .io_outer_finish_valid( L2BroadcastHub_io_outer_finish_valid ),
       .io_outer_finish_bits_header_src( L2BroadcastHub_io_outer_finish_bits_header_src ),
       .io_outer_finish_bits_header_dst( L2BroadcastHub_io_outer_finish_bits_header_dst ),
       .io_outer_finish_bits_payload_manager_xact_id( L2BroadcastHub_io_outer_finish_bits_payload_manager_xact_id ),
       .io_incoherent_1( io_incoherent_1 ),
       .io_incoherent_0( io_incoherent_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign L2BroadcastHub.io_outer_finish_ready = {1{$random}};
// synthesis translate_on
`endif
  TagCache tagCache(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( tagCache_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_uncached_acquire_bits_header_src( L2BroadcastHub_io_outer_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( L2BroadcastHub_io_outer_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( L2BroadcastHub_io_outer_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( L2BroadcastHub_io_outer_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_uncached( L2BroadcastHub_io_outer_acquire_bits_payload_uncached ),
       .io_uncached_acquire_bits_payload_a_type( L2BroadcastHub_io_outer_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_subblock( L2BroadcastHub_io_outer_acquire_bits_payload_subblock ),
       .io_uncached_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_uncached_grant_valid( tagCache_io_uncached_grant_valid ),
       .io_uncached_grant_bits_header_src( tagCache_io_uncached_grant_bits_header_src ),
       .io_uncached_grant_bits_header_dst( tagCache_io_uncached_grant_bits_header_dst ),
       .io_uncached_grant_bits_payload_data( tagCache_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( tagCache_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_manager_xact_id( tagCache_io_uncached_grant_bits_payload_manager_xact_id ),
       .io_uncached_grant_bits_payload_uncached( tagCache_io_uncached_grant_bits_payload_uncached ),
       .io_uncached_grant_bits_payload_g_type( tagCache_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( L2BroadcastHub_io_outer_finish_valid ),
       .io_uncached_finish_bits_header_src( L2BroadcastHub_io_outer_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( L2BroadcastHub_io_outer_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_manager_xact_id( L2BroadcastHub_io_outer_finish_bits_payload_manager_xact_id ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( tagCache_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( tagCache_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( tagCache_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( tagCache_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( tagCache_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( tagCache_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [135:0] io_enq_bits_payload_data,
    input  io_enq_bits_payload_uncached,
    input [1:0] io_enq_bits_payload_a_type,
    input [128:0] io_enq_bits_payload_subblock,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[135:0] io_deq_bits_payload_data,
    output io_deq_bits_payload_uncached,
    output[1:0] io_deq_bits_payload_a_type,
    output[128:0] io_deq_bits_payload_subblock,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[128:0] T10;
  wire[299:0] T11;
  reg [299:0] ram [1:0];
  wire[299:0] T12;
  wire[299:0] T13;
  wire[299:0] T14;
  wire[267:0] T15;
  wire[130:0] T16;
  wire[136:0] T17;
  wire[31:0] T18;
  wire[27:0] T19;
  wire[3:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[135:0] T23;
  wire[1:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {10{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_subblock = T10;
  assign T10 = T11[8'h80:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_a_type, io_enq_bits_payload_subblock};
  assign T17 = {io_enq_bits_payload_data, io_enq_bits_payload_uncached};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_a_type = T21;
  assign T21 = T11[8'h82:8'h81];
  assign io_deq_bits_payload_uncached = T22;
  assign T22 = T11[8'h83:8'h83];
  assign io_deq_bits_payload_data = T23;
  assign T23 = T11[9'h10b:8'h84];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T11[9'h10d:9'h10c];
  assign io_deq_bits_payload_addr = T25;
  assign T25 = T11[9'h127:9'h10e];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[9'h129:9'h128];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[9'h12b:9'h12a];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [135:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[135:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T27;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T28;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T29;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[170:0] T11;
  reg [170:0] ram [1:0];
  wire[170:0] T12;
  wire[170:0] T13;
  wire[170:0] T14;
  wire[140:0] T15;
  wire[138:0] T16;
  wire[29:0] T17;
  wire[27:0] T18;
  wire[135:0] T19;
  wire[1:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire empty;
  wire T25;
  wire T26;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T27 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T28 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T29 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_r_type = T10;
  assign T10 = T11[2'h2:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T17, T15};
  assign T15 = {io_enq_bits_payload_client_xact_id, T16};
  assign T16 = {io_enq_bits_payload_data, io_enq_bits_payload_r_type};
  assign T17 = {io_enq_bits_header_src, T18};
  assign T18 = {io_enq_bits_header_dst, io_enq_bits_payload_addr};
  assign io_deq_bits_payload_data = T19;
  assign T19 = T11[8'h8a:2'h3];
  assign io_deq_bits_payload_client_xact_id = T20;
  assign T20 = T11[8'h8c:8'h8b];
  assign io_deq_bits_payload_addr = T21;
  assign T21 = T11[8'ha6:8'h8d];
  assign io_deq_bits_header_dst = T22;
  assign T22 = T11[8'ha8:8'ha7];
  assign io_deq_bits_header_src = T23;
  assign T23 = T11[8'haa:8'ha9];
  assign io_deq_valid = T24;
  assign T24 = empty ^ 1'h1;
  assign empty = ptr_match & T25;
  assign T25 = maybe_full ^ 1'h1;
  assign io_enq_ready = T26;
  assign T26 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[7:0] T11;
  reg [7:0] ram [1:0];
  wire[7:0] T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[5:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_manager_xact_id = T10;
  assign T10 = T11[2'h3:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_header_src, T15};
  assign T15 = {io_enq_bits_header_dst, io_enq_bits_payload_manager_xact_id};
  assign io_deq_bits_header_dst = T16;
  assign T16 = T11[3'h5:3'h4];
  assign io_deq_bits_header_src = T17;
  assign T17 = T11[3'h7:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [135:0] io_enq_bits_payload_data,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [3:0] io_enq_bits_payload_manager_xact_id,
    input  io_enq_bits_payload_uncached,
    input [1:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[135:0] io_deq_bits_payload_data,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[3:0] io_deq_bits_payload_manager_xact_id,
    output io_deq_bits_payload_uncached,
    output[1:0] io_deq_bits_payload_g_type,
    output[2:0] io_count
);

  wire[2:0] T0;
  wire[1:0] ptr_diff;
  reg [1:0] R1;
  wire[1:0] T30;
  wire[1:0] T2;
  wire[1:0] T3;
  wire do_deq;
  reg [1:0] R4;
  wire[1:0] T31;
  wire[1:0] T5;
  wire[1:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T32;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[148:0] T11;
  reg [148:0] ram [3:0];
  wire[148:0] T12;
  wire[148:0] T13;
  wire[148:0] T14;
  wire[8:0] T15;
  wire[2:0] T16;
  wire[5:0] T17;
  wire[139:0] T18;
  wire[137:0] T19;
  wire T20;
  wire[3:0] T21;
  wire[1:0] T22;
  wire[135:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire T29;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T30 = reset ? 2'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 2'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T31 = reset ? 2'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 2'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T32 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_g_type = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_uncached, io_enq_bits_payload_g_type};
  assign T17 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_manager_xact_id};
  assign T18 = {io_enq_bits_header_src, T19};
  assign T19 = {io_enq_bits_header_dst, io_enq_bits_payload_data};
  assign io_deq_bits_payload_uncached = T20;
  assign T20 = T11[2'h2:2'h2];
  assign io_deq_bits_payload_manager_xact_id = T21;
  assign T21 = T11[3'h6:2'h3];
  assign io_deq_bits_payload_client_xact_id = T22;
  assign T22 = T11[4'h8:3'h7];
  assign io_deq_bits_payload_data = T23;
  assign T23 = T11[8'h90:4'h9];
  assign io_deq_bits_header_dst = T24;
  assign T24 = T11[8'h92:8'h91];
  assign io_deq_bits_header_src = T25;
  assign T25 = T11[8'h94:8'h93];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = T29 | io_deq_ready;
  assign T29 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 2'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 2'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_p_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T23;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T24;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[27:0] T15;
  wire[3:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_p_type = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_payload_addr, io_enq_bits_payload_p_type};
  assign T16 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_addr = T17;
  assign T17 = T11[5'h1b:2'h2];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T11[5'h1d:5'h1c];
  assign io_deq_bits_header_src = T19;
  assign T19 = T11[5'h1f:5'h1e];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [135:0] io_tiles_0_acquire_bits_payload_data,
    input  io_tiles_0_acquire_bits_payload_uncached,
    input [1:0] io_tiles_0_acquire_bits_payload_a_type,
    input [128:0] io_tiles_0_acquire_bits_payload_subblock,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[135:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_manager_xact_id,
    output io_tiles_0_grant_bits_payload_uncached,
    output[1:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [3:0] io_tiles_0_finish_bits_payload_manager_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [135:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[4:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr,
    input  io_incoherent_0
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire[3:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[135:0] T5;
  wire[1:0] T6;
  wire[25:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire[128:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[135:0] T14;
  wire[1:0] T15;
  wire[25:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire[3:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[135:0] T25;
  wire[1:0] T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire[128:0] T31;
  wire[1:0] T32;
  wire T33;
  wire[135:0] T34;
  wire[1:0] T35;
  wire[25:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_pcr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire[4:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_payload_addr;
  wire[1:0] htif_io_mem_acquire_bits_payload_client_xact_id;
  wire[135:0] htif_io_mem_acquire_bits_payload_data;
  wire htif_io_mem_acquire_bits_payload_uncached;
  wire[1:0] htif_io_mem_acquire_bits_payload_a_type;
  wire[128:0] htif_io_mem_acquire_bits_payload_subblock;
  wire htif_io_mem_grant_ready;
  wire htif_io_mem_finish_valid;
  wire[1:0] htif_io_mem_finish_bits_header_dst;
  wire[3:0] htif_io_mem_finish_bits_payload_manager_xact_id;
  wire htif_io_mem_probe_ready;
  wire htif_io_mem_release_valid;
  wire[25:0] htif_io_mem_release_bits_payload_addr;
  wire[1:0] htif_io_mem_release_bits_payload_client_xact_id;
  wire[135:0] htif_io_mem_release_bits_payload_data;
  wire[2:0] htif_io_mem_release_bits_payload_r_type;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[25:0] Queue_4_io_deq_bits_payload_addr;
  wire[1:0] Queue_4_io_deq_bits_payload_client_xact_id;
  wire[135:0] Queue_4_io_deq_bits_payload_data;
  wire Queue_4_io_deq_bits_payload_uncached;
  wire[1:0] Queue_4_io_deq_bits_payload_a_type;
  wire[128:0] Queue_4_io_deq_bits_payload_subblock;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[1:0] Queue_5_io_deq_bits_header_src;
  wire[1:0] Queue_5_io_deq_bits_header_dst;
  wire[25:0] Queue_5_io_deq_bits_payload_addr;
  wire[1:0] Queue_5_io_deq_bits_payload_client_xact_id;
  wire[135:0] Queue_5_io_deq_bits_payload_data;
  wire[2:0] Queue_5_io_deq_bits_payload_r_type;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[1:0] Queue_6_io_deq_bits_header_src;
  wire[1:0] Queue_6_io_deq_bits_header_dst;
  wire[3:0] Queue_6_io_deq_bits_payload_manager_xact_id;
  wire Queue_7_io_enq_ready;
  wire Queue_7_io_deq_valid;
  wire[1:0] Queue_7_io_deq_bits_header_src;
  wire[1:0] Queue_7_io_deq_bits_header_dst;
  wire[135:0] Queue_7_io_deq_bits_payload_data;
  wire[1:0] Queue_7_io_deq_bits_payload_client_xact_id;
  wire[3:0] Queue_7_io_deq_bits_payload_manager_xact_id;
  wire Queue_7_io_deq_bits_payload_uncached;
  wire[1:0] Queue_7_io_deq_bits_payload_g_type;
  wire Queue_8_io_enq_ready;
  wire Queue_8_io_deq_valid;
  wire[1:0] Queue_8_io_deq_bits_header_src;
  wire[1:0] Queue_8_io_deq_bits_header_dst;
  wire[25:0] Queue_8_io_deq_bits_payload_addr;
  wire[1:0] Queue_8_io_deq_bits_payload_p_type;
  wire Queue_9_io_enq_ready;
  wire Queue_9_io_deq_valid;
  wire[1:0] Queue_9_io_deq_bits_header_src;
  wire[1:0] Queue_9_io_deq_bits_header_dst;
  wire[25:0] Queue_9_io_deq_bits_payload_addr;
  wire[1:0] Queue_9_io_deq_bits_payload_client_xact_id;
  wire[135:0] Queue_9_io_deq_bits_payload_data;
  wire Queue_9_io_deq_bits_payload_uncached;
  wire[1:0] Queue_9_io_deq_bits_payload_a_type;
  wire[128:0] Queue_9_io_deq_bits_payload_subblock;
  wire Queue_10_io_enq_ready;
  wire Queue_10_io_deq_valid;
  wire[1:0] Queue_10_io_deq_bits_header_src;
  wire[1:0] Queue_10_io_deq_bits_header_dst;
  wire[25:0] Queue_10_io_deq_bits_payload_addr;
  wire[1:0] Queue_10_io_deq_bits_payload_client_xact_id;
  wire[135:0] Queue_10_io_deq_bits_payload_data;
  wire[2:0] Queue_10_io_deq_bits_payload_r_type;
  wire Queue_11_io_enq_ready;
  wire Queue_11_io_deq_valid;
  wire[1:0] Queue_11_io_deq_bits_header_src;
  wire[1:0] Queue_11_io_deq_bits_header_dst;
  wire[3:0] Queue_11_io_deq_bits_payload_manager_xact_id;
  wire Queue_12_io_enq_ready;
  wire Queue_12_io_deq_valid;
  wire[1:0] Queue_12_io_deq_bits_header_src;
  wire[1:0] Queue_12_io_deq_bits_header_dst;
  wire[135:0] Queue_12_io_deq_bits_payload_data;
  wire[1:0] Queue_12_io_deq_bits_payload_client_xact_id;
  wire[3:0] Queue_12_io_deq_bits_payload_manager_xact_id;
  wire Queue_12_io_deq_bits_payload_uncached;
  wire[1:0] Queue_12_io_deq_bits_payload_g_type;
  wire Queue_13_io_enq_ready;
  wire Queue_13_io_deq_valid;
  wire[1:0] Queue_13_io_deq_bits_header_src;
  wire[1:0] Queue_13_io_deq_bits_header_dst;
  wire[25:0] Queue_13_io_deq_bits_payload_addr;
  wire[1:0] Queue_13_io_deq_bits_payload_p_type;
  wire outmemsys_io_tiles_0_acquire_ready;
  wire outmemsys_io_tiles_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_dst;
  wire[135:0] outmemsys_io_tiles_0_grant_bits_payload_data;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_manager_xact_id;
  wire outmemsys_io_tiles_0_grant_bits_payload_uncached;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_payload_g_type;
  wire outmemsys_io_tiles_0_finish_ready;
  wire outmemsys_io_tiles_0_probe_valid;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_dst;
  wire[25:0] outmemsys_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_payload_p_type;
  wire outmemsys_io_tiles_0_release_ready;
  wire outmemsys_io_htif_acquire_ready;
  wire outmemsys_io_htif_grant_valid;
  wire[1:0] outmemsys_io_htif_grant_bits_header_src;
  wire[1:0] outmemsys_io_htif_grant_bits_header_dst;
  wire[135:0] outmemsys_io_htif_grant_bits_payload_data;
  wire[1:0] outmemsys_io_htif_grant_bits_payload_client_xact_id;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_manager_xact_id;
  wire outmemsys_io_htif_grant_bits_payload_uncached;
  wire[1:0] outmemsys_io_htif_grant_bits_payload_g_type;
  wire outmemsys_io_htif_finish_ready;
  wire outmemsys_io_htif_probe_valid;
  wire[1:0] outmemsys_io_htif_probe_bits_header_src;
  wire[1:0] outmemsys_io_htif_probe_bits_header_dst;
  wire[25:0] outmemsys_io_htif_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_htif_probe_bits_payload_p_type;
  wire outmemsys_io_htif_release_ready;
  wire outmemsys_io_mem_req_cmd_valid;
  wire[25:0] outmemsys_io_mem_req_cmd_bits_addr;
  wire[4:0] outmemsys_io_mem_req_cmd_bits_tag;
  wire outmemsys_io_mem_req_cmd_bits_rw;
  wire outmemsys_io_mem_req_data_valid;
  wire[127:0] outmemsys_io_mem_req_data_bits_data;


  assign T0 = htif_io_mem_finish_bits_payload_manager_xact_id;
  assign T1 = htif_io_mem_finish_bits_header_dst;
  assign T2 = 2'h1;
  assign T3 = htif_io_mem_finish_valid;
  assign T4 = htif_io_mem_release_bits_payload_r_type;
  assign T5 = htif_io_mem_release_bits_payload_data;
  assign T6 = htif_io_mem_release_bits_payload_client_xact_id;
  assign T7 = htif_io_mem_release_bits_payload_addr;
  assign T8 = 2'h0;
  assign T9 = 2'h1;
  assign T10 = htif_io_mem_release_valid;
  assign T11 = htif_io_mem_acquire_bits_payload_subblock;
  assign T12 = htif_io_mem_acquire_bits_payload_a_type;
  assign T13 = htif_io_mem_acquire_bits_payload_uncached;
  assign T14 = htif_io_mem_acquire_bits_payload_data;
  assign T15 = htif_io_mem_acquire_bits_payload_client_xact_id;
  assign T16 = htif_io_mem_acquire_bits_payload_addr;
  assign T17 = 2'h0;
  assign T18 = 2'h1;
  assign T19 = htif_io_mem_acquire_valid;
  assign T20 = io_tiles_0_finish_bits_payload_manager_xact_id;
  assign T21 = io_tiles_0_finish_bits_header_dst;
  assign T22 = 2'h0;
  assign T23 = io_tiles_0_finish_valid;
  assign T24 = io_tiles_0_release_bits_payload_r_type;
  assign T25 = io_tiles_0_release_bits_payload_data;
  assign T26 = io_tiles_0_release_bits_payload_client_xact_id;
  assign T27 = io_tiles_0_release_bits_payload_addr;
  assign T28 = 2'h0;
  assign T29 = 2'h0;
  assign T30 = io_tiles_0_release_valid;
  assign T31 = io_tiles_0_acquire_bits_payload_subblock;
  assign T32 = io_tiles_0_acquire_bits_payload_a_type;
  assign T33 = io_tiles_0_acquire_bits_payload_uncached;
  assign T34 = io_tiles_0_acquire_bits_payload_data;
  assign T35 = io_tiles_0_acquire_bits_payload_client_xact_id;
  assign T36 = io_tiles_0_acquire_bits_payload_addr;
  assign T37 = 2'h0;
  assign T38 = 2'h0;
  assign T39 = io_tiles_0_acquire_valid;
  assign T40 = Queue_10_io_enq_ready;
  assign T41 = Queue_11_io_enq_ready;
  assign T42 = Queue_9_io_enq_ready;
//  assign io_mem_backup_req_bits = {1{$random}};
//  assign io_mem_backup_req_valid = {1{$random}};
  assign io_htif_0_ipi_rep_bits = {1{$random}};
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
//  assign io_htif_0_id = {1{$random}};
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_tiles_0_release_ready = T43;
  assign T43 = Queue_5_io_enq_ready;
  assign io_tiles_0_probe_bits_payload_p_type = Queue_8_io_deq_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_addr = Queue_8_io_deq_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = Queue_8_io_deq_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = Queue_8_io_deq_bits_header_src;
  assign io_tiles_0_probe_valid = Queue_8_io_deq_valid;
  assign io_tiles_0_finish_ready = T44;
  assign T44 = Queue_6_io_enq_ready;
  assign io_tiles_0_grant_bits_payload_g_type = Queue_7_io_deq_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_uncached = Queue_7_io_deq_bits_payload_uncached;
  assign io_tiles_0_grant_bits_payload_manager_xact_id = Queue_7_io_deq_bits_payload_manager_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = Queue_7_io_deq_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = Queue_7_io_deq_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = Queue_7_io_deq_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = Queue_7_io_deq_bits_header_src;
  assign io_tiles_0_grant_valid = Queue_7_io_deq_valid;
  assign io_tiles_0_acquire_ready = T45;
  assign T45 = Queue_4_io_enq_ready;
//  assign io_mem_resp_ready = {1{$random}};
  assign io_mem_req_data_bits_data = outmemsys_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = outmemsys_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = outmemsys_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = outmemsys_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = outmemsys_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = outmemsys_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = htif_io_host_debug_stats_pcr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_pcr( htif_io_host_debug_stats_pcr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( T42 ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( htif_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( htif_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( htif_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_uncached( htif_io_mem_acquire_bits_payload_uncached ),
       .io_mem_acquire_bits_payload_a_type( htif_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_subblock( htif_io_mem_acquire_bits_payload_subblock ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( Queue_12_io_deq_valid ),
       .io_mem_grant_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_mem_grant_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_mem_grant_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_manager_xact_id( Queue_12_io_deq_bits_payload_manager_xact_id ),
       .io_mem_grant_bits_payload_uncached( Queue_12_io_deq_bits_payload_uncached ),
       .io_mem_grant_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type ),
       .io_mem_finish_ready( T41 ),
       .io_mem_finish_valid( htif_io_mem_finish_valid ),
       //.io_mem_finish_bits_header_src(  )
       .io_mem_finish_bits_header_dst( htif_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_manager_xact_id( htif_io_mem_finish_bits_payload_manager_xact_id ),
       .io_mem_probe_ready( htif_io_mem_probe_ready ),
       .io_mem_probe_valid( Queue_13_io_deq_valid ),
       .io_mem_probe_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_mem_probe_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_mem_probe_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type ),
       .io_mem_release_ready( T40 ),
       .io_mem_release_valid( htif_io_mem_release_valid ),
       //.io_mem_release_bits_header_src(  )
       //.io_mem_release_bits_header_dst(  )
       .io_mem_release_bits_payload_addr( htif_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( htif_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_data( htif_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( htif_io_mem_release_bits_payload_r_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign htif.io_mem_release_bits_payload_addr = {1{$random}};
    assign htif.io_mem_release_bits_payload_client_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_data = {5{$random}};
    assign htif.io_mem_release_bits_payload_r_type = {1{$random}};
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
// synthesis translate_on
`endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_0_acquire_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Queue_4_io_deq_valid ),
       .io_tiles_0_acquire_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_uncached( Queue_4_io_deq_bits_payload_uncached ),
       .io_tiles_0_acquire_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_subblock( Queue_4_io_deq_bits_payload_subblock ),
       .io_tiles_0_grant_ready( Queue_7_io_enq_ready ),
       .io_tiles_0_grant_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_manager_xact_id( outmemsys_io_tiles_0_grant_bits_payload_manager_xact_id ),
       .io_tiles_0_grant_bits_payload_uncached( outmemsys_io_tiles_0_grant_bits_payload_uncached ),
       .io_tiles_0_grant_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Queue_6_io_deq_valid ),
       .io_tiles_0_finish_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_manager_xact_id( Queue_6_io_deq_bits_payload_manager_xact_id ),
       .io_tiles_0_probe_ready( Queue_8_io_enq_ready ),
       .io_tiles_0_probe_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( outmemsys_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Queue_5_io_deq_valid ),
       .io_tiles_0_release_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type ),
       .io_htif_acquire_ready( outmemsys_io_htif_acquire_ready ),
       .io_htif_acquire_valid( Queue_9_io_deq_valid ),
       .io_htif_acquire_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_htif_acquire_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_htif_acquire_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_htif_acquire_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_htif_acquire_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_htif_acquire_bits_payload_uncached( Queue_9_io_deq_bits_payload_uncached ),
       .io_htif_acquire_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_htif_acquire_bits_payload_subblock( Queue_9_io_deq_bits_payload_subblock ),
       .io_htif_grant_ready( Queue_12_io_enq_ready ),
       .io_htif_grant_valid( outmemsys_io_htif_grant_valid ),
       .io_htif_grant_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_htif_grant_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_htif_grant_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_htif_grant_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_htif_grant_bits_payload_manager_xact_id( outmemsys_io_htif_grant_bits_payload_manager_xact_id ),
       .io_htif_grant_bits_payload_uncached( outmemsys_io_htif_grant_bits_payload_uncached ),
       .io_htif_grant_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_htif_finish_ready( outmemsys_io_htif_finish_ready ),
       .io_htif_finish_valid( Queue_11_io_deq_valid ),
       .io_htif_finish_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_htif_finish_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_htif_finish_bits_payload_manager_xact_id( Queue_11_io_deq_bits_payload_manager_xact_id ),
       .io_htif_probe_ready( Queue_13_io_enq_ready ),
       .io_htif_probe_valid( outmemsys_io_htif_probe_valid ),
       .io_htif_probe_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_htif_probe_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_htif_probe_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_htif_probe_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_htif_release_ready( outmemsys_io_htif_release_ready ),
       .io_htif_release_valid( Queue_10_io_deq_valid ),
       .io_htif_release_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_htif_release_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_htif_release_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_htif_release_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_htif_release_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_htif_release_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type ),
       .io_incoherent_1( 1'h1 ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( outmemsys_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( outmemsys_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( outmemsys_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( outmemsys_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( outmemsys_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( outmemsys_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( T39 ),
       .io_enq_bits_header_src( T38 ),
       .io_enq_bits_header_dst( T37 ),
       .io_enq_bits_payload_addr( T36 ),
       .io_enq_bits_payload_client_xact_id( T35 ),
       .io_enq_bits_payload_data( T34 ),
       .io_enq_bits_payload_uncached( T33 ),
       .io_enq_bits_payload_a_type( T32 ),
       .io_enq_bits_payload_subblock( T31 ),
       .io_deq_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_deq_bits_payload_uncached( Queue_4_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_subblock( Queue_4_io_deq_bits_payload_subblock )
       //.io_count(  )
  );
  Queue_4 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( T30 ),
       .io_enq_bits_header_src( T29 ),
       .io_enq_bits_header_dst( T28 ),
       .io_enq_bits_payload_addr( T27 ),
       .io_enq_bits_payload_client_xact_id( T26 ),
       .io_enq_bits_payload_data( T25 ),
       .io_enq_bits_payload_r_type( T24 ),
       .io_deq_ready( outmemsys_io_tiles_0_release_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type )
       //.io_count(  )
  );
  Queue_5 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( T23 ),
       .io_enq_bits_header_src( T22 ),
       .io_enq_bits_header_dst( T21 ),
       .io_enq_bits_payload_manager_xact_id( T20 ),
       .io_deq_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( Queue_6_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
  Queue_6 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_manager_xact_id( outmemsys_io_tiles_0_grant_bits_payload_manager_xact_id ),
       .io_enq_bits_payload_uncached( outmemsys_io_tiles_0_grant_bits_payload_uncached ),
       .io_enq_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_deq_ready( io_tiles_0_grant_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_7_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_7_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_manager_xact_id( Queue_7_io_deq_bits_payload_manager_xact_id ),
       .io_deq_bits_payload_uncached( Queue_7_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_g_type( Queue_7_io_deq_bits_payload_g_type )
       //.io_count(  )
  );
  Queue_7 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_enq_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_deq_ready( io_tiles_0_probe_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_8_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_p_type( Queue_8_io_deq_bits_payload_p_type )
       //.io_count(  )
  );
  Queue_3 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( T19 ),
       .io_enq_bits_header_src( T18 ),
       .io_enq_bits_header_dst( T17 ),
       .io_enq_bits_payload_addr( T16 ),
       .io_enq_bits_payload_client_xact_id( T15 ),
       .io_enq_bits_payload_data( T14 ),
       .io_enq_bits_payload_uncached( T13 ),
       .io_enq_bits_payload_a_type( T12 ),
       .io_enq_bits_payload_subblock( T11 ),
       .io_deq_ready( outmemsys_io_htif_acquire_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_deq_bits_payload_uncached( Queue_9_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_subblock( Queue_9_io_deq_bits_payload_subblock )
       //.io_count(  )
  );
  Queue_4 Queue_10(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_10_io_enq_ready ),
       .io_enq_valid( T10 ),
       .io_enq_bits_header_src( T9 ),
       .io_enq_bits_header_dst( T8 ),
       .io_enq_bits_payload_addr( T7 ),
       .io_enq_bits_payload_client_xact_id( T6 ),
       .io_enq_bits_payload_data( T5 ),
       .io_enq_bits_payload_r_type( T4 ),
       .io_deq_ready( outmemsys_io_htif_release_ready ),
       .io_deq_valid( Queue_10_io_deq_valid ),
       .io_deq_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type )
       //.io_count(  )
  );
  Queue_5 Queue_11(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_11_io_enq_ready ),
       .io_enq_valid( T3 ),
       .io_enq_bits_header_src( T2 ),
       .io_enq_bits_header_dst( T1 ),
       .io_enq_bits_payload_manager_xact_id( T0 ),
       .io_deq_ready( outmemsys_io_htif_finish_ready ),
       .io_deq_valid( Queue_11_io_deq_valid ),
       .io_deq_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( Queue_11_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
  Queue_6 Queue_12(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_12_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_manager_xact_id( outmemsys_io_htif_grant_bits_payload_manager_xact_id ),
       .io_enq_bits_payload_uncached( outmemsys_io_htif_grant_bits_payload_uncached ),
       .io_enq_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_deq_ready( htif_io_mem_grant_ready ),
       .io_deq_valid( Queue_12_io_deq_valid ),
       .io_deq_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_manager_xact_id( Queue_12_io_deq_bits_payload_manager_xact_id ),
       .io_deq_bits_payload_uncached( Queue_12_io_deq_bits_payload_uncached ),
       .io_deq_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type )
       //.io_count(  )
  );
  Queue_7 Queue_13(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_13_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_enq_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_deq_ready( htif_io_mem_probe_ready ),
       .io_deq_valid( Queue_13_io_deq_valid ),
       .io_deq_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type )
       //.io_count(  )
  );
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [4:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[4:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[69:0] T11;
  reg [69:0] ram [1:0];
  wire[69:0] T12;
  wire[69:0] T13;
  wire[69:0] T14;
  wire[68:0] T15;
  wire[4:0] T16;
  wire T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_rw, T15};
  assign T15 = {io_enq_bits_addr, io_enq_bits_data};
  assign io_deq_bits_addr = T16;
  assign T16 = T11[7'h44:7'h40];
  assign io_deq_bits_rw = T17;
  assign T17 = T11[7'h45:7'h45];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[63:0] T10;
  reg [63:0] ram [1:0];
  wire[63:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire T10;
  reg [0:0] ram [1:0];
  wire T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    input  io_mem_backup_en,
    output io_in_mem_ready,
    input  io_in_mem_valid,
    input  io_out_mem_ready,
    output io_out_mem_valid
);

  wire resetSigs_0;
  reg  R0;
  reg  R1;
  wire Queue_0_io_enq_ready;
  wire Queue_0_io_deq_valid;
  wire Queue_0_io_deq_bits_rw;
  wire[4:0] Queue_0_io_deq_bits_addr;
  wire[63:0] Queue_0_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire Queue_2_io_deq_bits;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire Queue_3_io_deq_bits;
  wire RocketTile_io_tilelink_acquire_valid;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_header_src;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_header_dst;
  wire[25:0] RocketTile_io_tilelink_acquire_bits_payload_addr;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_payload_client_xact_id;
  wire[135:0] RocketTile_io_tilelink_acquire_bits_payload_data;
  wire RocketTile_io_tilelink_acquire_bits_payload_uncached;
  wire[1:0] RocketTile_io_tilelink_acquire_bits_payload_a_type;
  wire[128:0] RocketTile_io_tilelink_acquire_bits_payload_subblock;
  wire RocketTile_io_tilelink_grant_ready;
  wire RocketTile_io_tilelink_finish_valid;
  wire[1:0] RocketTile_io_tilelink_finish_bits_header_src;
  wire[1:0] RocketTile_io_tilelink_finish_bits_header_dst;
  wire[3:0] RocketTile_io_tilelink_finish_bits_payload_manager_xact_id;
  wire RocketTile_io_tilelink_probe_ready;
  wire RocketTile_io_tilelink_release_valid;
  wire[1:0] RocketTile_io_tilelink_release_bits_header_src;
  wire[1:0] RocketTile_io_tilelink_release_bits_header_dst;
  wire[25:0] RocketTile_io_tilelink_release_bits_payload_addr;
  wire[1:0] RocketTile_io_tilelink_release_bits_payload_client_xact_id;
  wire[135:0] RocketTile_io_tilelink_release_bits_payload_data;
  wire[2:0] RocketTile_io_tilelink_release_bits_payload_r_type;
  wire RocketTile_io_host_pcr_req_ready;
  wire RocketTile_io_host_pcr_rep_valid;
  wire[63:0] RocketTile_io_host_pcr_rep_bits;
  wire RocketTile_io_host_ipi_req_valid;
  wire RocketTile_io_host_ipi_req_bits;
  wire RocketTile_io_host_ipi_rep_ready;
  wire RocketTile_io_host_debug_stats_pcr;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_pcr;
  wire uncore_io_mem_req_cmd_valid;
  wire[25:0] uncore_io_mem_req_cmd_bits_addr;
  wire[4:0] uncore_io_mem_req_cmd_bits_tag;
  wire uncore_io_mem_req_cmd_bits_rw;
  wire uncore_io_mem_req_data_valid;
  wire[127:0] uncore_io_mem_req_data_bits_data;
  wire uncore_io_tiles_0_acquire_ready;
  wire uncore_io_tiles_0_grant_valid;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_src;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_dst;
  wire[135:0] uncore_io_tiles_0_grant_bits_payload_data;
  wire[1:0] uncore_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_manager_xact_id;
  wire uncore_io_tiles_0_grant_bits_payload_uncached;
  wire[1:0] uncore_io_tiles_0_grant_bits_payload_g_type;
  wire uncore_io_tiles_0_finish_ready;
  wire uncore_io_tiles_0_probe_valid;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_src;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_dst;
  wire[25:0] uncore_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] uncore_io_tiles_0_probe_bits_payload_p_type;
  wire uncore_io_tiles_0_release_ready;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_pcr_req_valid;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire[4:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire uncore_io_htif_0_ipi_req_ready;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_rep_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign resetSigs_0 = uncore_io_htif_0_reset;
//  assign io_out_mem_valid = {1{$random}};
//  assign io_in_mem_ready = {1{$random}};
//  assign io_mem_resp_ready = {1{$random}};
  assign io_mem_req_data_bits_data = uncore_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = uncore_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = uncore_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = uncore_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = uncore_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = uncore_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = uncore_io_host_debug_stats_pcr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
  RocketTile RocketTile(.clk(clk), .reset(resetSigs_0),
       .io_tilelink_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tilelink_acquire_valid( RocketTile_io_tilelink_acquire_valid ),
       .io_tilelink_acquire_bits_header_src( RocketTile_io_tilelink_acquire_bits_header_src ),
       .io_tilelink_acquire_bits_header_dst( RocketTile_io_tilelink_acquire_bits_header_dst ),
       .io_tilelink_acquire_bits_payload_addr( RocketTile_io_tilelink_acquire_bits_payload_addr ),
       .io_tilelink_acquire_bits_payload_client_xact_id( RocketTile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tilelink_acquire_bits_payload_data( RocketTile_io_tilelink_acquire_bits_payload_data ),
       .io_tilelink_acquire_bits_payload_uncached( RocketTile_io_tilelink_acquire_bits_payload_uncached ),
       .io_tilelink_acquire_bits_payload_a_type( RocketTile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tilelink_acquire_bits_payload_subblock( RocketTile_io_tilelink_acquire_bits_payload_subblock ),
       .io_tilelink_grant_ready( RocketTile_io_tilelink_grant_ready ),
       .io_tilelink_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tilelink_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tilelink_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tilelink_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tilelink_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tilelink_grant_bits_payload_manager_xact_id( uncore_io_tiles_0_grant_bits_payload_manager_xact_id ),
       .io_tilelink_grant_bits_payload_uncached( uncore_io_tiles_0_grant_bits_payload_uncached ),
       .io_tilelink_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tilelink_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tilelink_finish_valid( RocketTile_io_tilelink_finish_valid ),
       .io_tilelink_finish_bits_header_src( RocketTile_io_tilelink_finish_bits_header_src ),
       .io_tilelink_finish_bits_header_dst( RocketTile_io_tilelink_finish_bits_header_dst ),
       .io_tilelink_finish_bits_payload_manager_xact_id( RocketTile_io_tilelink_finish_bits_payload_manager_xact_id ),
       .io_tilelink_probe_ready( RocketTile_io_tilelink_probe_ready ),
       .io_tilelink_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tilelink_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tilelink_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tilelink_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tilelink_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tilelink_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tilelink_release_valid( RocketTile_io_tilelink_release_valid ),
       .io_tilelink_release_bits_header_src( RocketTile_io_tilelink_release_bits_header_src ),
       .io_tilelink_release_bits_header_dst( RocketTile_io_tilelink_release_bits_header_dst ),
       .io_tilelink_release_bits_payload_addr( RocketTile_io_tilelink_release_bits_payload_addr ),
       .io_tilelink_release_bits_payload_client_xact_id( RocketTile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tilelink_release_bits_payload_data( RocketTile_io_tilelink_release_bits_payload_data ),
       .io_tilelink_release_bits_payload_r_type( RocketTile_io_tilelink_release_bits_payload_r_type ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( RocketTile_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_0_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_0_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( RocketTile_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( RocketTile_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( RocketTile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( RocketTile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_pcr( RocketTile_io_host_debug_stats_pcr )
  );
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_pcr( uncore_io_host_debug_stats_pcr ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( uncore_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( uncore_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( uncore_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( uncore_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( uncore_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( uncore_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_tiles_0_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( RocketTile_io_tilelink_acquire_valid ),
       .io_tiles_0_acquire_bits_header_src( RocketTile_io_tilelink_acquire_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( RocketTile_io_tilelink_acquire_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( RocketTile_io_tilelink_acquire_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( RocketTile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( RocketTile_io_tilelink_acquire_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_uncached( RocketTile_io_tilelink_acquire_bits_payload_uncached ),
       .io_tiles_0_acquire_bits_payload_a_type( RocketTile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_subblock( RocketTile_io_tilelink_acquire_bits_payload_subblock ),
       .io_tiles_0_grant_ready( RocketTile_io_tilelink_grant_ready ),
       .io_tiles_0_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_manager_xact_id( uncore_io_tiles_0_grant_bits_payload_manager_xact_id ),
       .io_tiles_0_grant_bits_payload_uncached( uncore_io_tiles_0_grant_bits_payload_uncached ),
       .io_tiles_0_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( RocketTile_io_tilelink_finish_valid ),
       .io_tiles_0_finish_bits_header_src( RocketTile_io_tilelink_finish_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( RocketTile_io_tilelink_finish_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_manager_xact_id( RocketTile_io_tilelink_finish_bits_payload_manager_xact_id ),
       .io_tiles_0_probe_ready( RocketTile_io_tilelink_probe_ready ),
       .io_tiles_0_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( RocketTile_io_tilelink_release_valid ),
       .io_tiles_0_release_bits_header_src( RocketTile_io_tilelink_release_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( RocketTile_io_tilelink_release_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( RocketTile_io_tilelink_release_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( RocketTile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_data( RocketTile_io_tilelink_release_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( RocketTile_io_tilelink_release_bits_payload_r_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_0_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_pcr( RocketTile_io_host_debug_stats_pcr ),
       .io_incoherent_0( uncore_io_htif_0_reset )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
// synthesis translate_on
`endif
  Queue_0 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( RocketTile_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_0_io_deq_bits_data )
       //.io_count(  )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_pcr_rep_valid ),
       .io_enq_bits( RocketTile_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_ipi_req_valid ),
       .io_enq_bits( RocketTile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module DataArray_T6(
  input CLK,
  input RST,
  input init,
  input [8:0] W0A,
  input W0E,
  input [135:0] W0I,
  input [135:0] W0M,
  input [8:0] R1A,
  input R1E,
  output [135:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+68) begin
    for (j=1; j<68; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [135:0] ram [511:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {5 {$random}};
    end
  `endif
  reg [8:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][67:0] <= W0I[67:0];
  if (W0E && W0M[68]) ram[W0A][135:68] <= W0I[135:68];
end
assign R1O = ram[reg_R1A];

endmodule


module TagCacheDataArray_T2(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0M,
  input [127:0] RW0I,
  output [127:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<4; i=i+32) begin
    for (j=1; j<32; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][31:0] <= RW0I[31:0];
  if (RW0E && RW0W && RW0M[32]) ram[RW0A][63:32] <= RW0I[63:32];
  if (RW0E && RW0W && RW0M[64]) ram[RW0A][95:64] <= RW0I[95:64];
  if (RW0E && RW0W && RW0M[96]) ram[RW0A][127:96] <= RW0I[127:96];
end
assign RW0O = ram[reg_RW0A];

endmodule


module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [6:0] W0A,
  input W0E,
  input [83:0] W0I,
  input [83:0] W0M,
  input [6:0] R1A,
  input R1E,
  output [83:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<4; i=i+21) begin
    for (j=1; j<21; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [83:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
    end
  `endif
  reg [6:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][20:0] <= W0I[20:0];
  if (W0E && W0M[21]) ram[W0A][41:21] <= W0I[41:21];
  if (W0E && W0M[42]) ram[W0A][62:42] <= W0I[62:42];
  if (W0E && W0M[63]) ram[W0A][83:63] <= W0I[83:63];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [6:0] RW0A,
  input RW0E,
  input RW0W,
  input [37:0] RW0M,
  input [37:0] RW0I,
  output [37:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+19) begin
    for (j=1; j<19; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [37:0] ram [127:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {2 {$random}};
    end
  `endif
  reg [6:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][18:0] <= RW0I[18:0];
  if (RW0E && RW0W && RW0M[19]) ram[RW0A][37:19] <= RW0I[37:19];
end
assign RW0O = ram[reg_RW0A];

endmodule


module TagCacheMetadataArray_metaArray(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [135:0] W0I,
  input [135:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [135:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<8; i=i+17) begin
    for (j=1; j<17; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [135:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {5 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][16:0] <= W0I[16:0];
  if (W0E && W0M[17]) ram[W0A][33:17] <= W0I[33:17];
  if (W0E && W0M[34]) ram[W0A][50:34] <= W0I[50:34];
  if (W0E && W0M[51]) ram[W0A][67:51] <= W0I[67:51];
  if (W0E && W0M[68]) ram[W0A][84:68] <= W0I[84:68];
  if (W0E && W0M[85]) ram[W0A][101:85] <= W0I[101:85];
  if (W0E && W0M[102]) ram[W0A][118:102] <= W0I[118:102];
  if (W0E && W0M[119]) ram[W0A][135:119] <= W0I[135:119];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_T168(
  input CLK,
  input RST,
  input init,
  input [8:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [511:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [8:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


